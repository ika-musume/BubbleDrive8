module PositionPageConverter 
(
    input   wire            nCONV,
    input   wire    [11:0]  POS,
    output  reg     [11:0]  PAGE = 12'd4095
);

    always @ (negedge nCONV)
    begin
        case (POS)
            12'd0: PAGE <= 12'd1862;
            12'd1: PAGE <= 12'd331;
            12'd2: PAGE <= 12'd853;
            12'd3: PAGE <= 12'd1375;
            12'd4: PAGE <= 12'd1897;
            12'd5: PAGE <= 12'd366;
            12'd6: PAGE <= 12'd888;
            12'd7: PAGE <= 12'd1410;
            12'd8: PAGE <= 12'd1932;
            12'd9: PAGE <= 12'd401;
            12'd10: PAGE <= 12'd923;
            12'd11: PAGE <= 12'd1445;
            12'd12: PAGE <= 12'd1967;
            12'd13: PAGE <= 12'd436;
            12'd14: PAGE <= 12'd958;
            12'd15: PAGE <= 12'd1480;
            12'd16: PAGE <= 12'd2002;
            12'd17: PAGE <= 12'd471;
            12'd18: PAGE <= 12'd993;
            12'd19: PAGE <= 12'd1515;
            12'd20: PAGE <= 12'd2037;
            12'd21: PAGE <= 12'd506;
            12'd22: PAGE <= 12'd1028;
            12'd23: PAGE <= 12'd1550;
            12'd24: PAGE <= 12'd19;
            12'd25: PAGE <= 12'd541;
            12'd26: PAGE <= 12'd1063;
            12'd27: PAGE <= 12'd1585;
            12'd28: PAGE <= 12'd54;
            12'd29: PAGE <= 12'd576;
            12'd30: PAGE <= 12'd1098;
            12'd31: PAGE <= 12'd1620;
            12'd32: PAGE <= 12'd89;
            12'd33: PAGE <= 12'd611;
            12'd34: PAGE <= 12'd1133;
            12'd35: PAGE <= 12'd1655;
            12'd36: PAGE <= 12'd124;
            12'd37: PAGE <= 12'd646;
            12'd38: PAGE <= 12'd1168;
            12'd39: PAGE <= 12'd1690;
            12'd40: PAGE <= 12'd159;
            12'd41: PAGE <= 12'd681;
            12'd42: PAGE <= 12'd1203;
            12'd43: PAGE <= 12'd1725;
            12'd44: PAGE <= 12'd194;
            12'd45: PAGE <= 12'd716;
            12'd46: PAGE <= 12'd1238;
            12'd47: PAGE <= 12'd1760;
            12'd48: PAGE <= 12'd229;
            12'd49: PAGE <= 12'd751;
            12'd50: PAGE <= 12'd1273;
            12'd51: PAGE <= 12'd1795;
            12'd52: PAGE <= 12'd264;
            12'd53: PAGE <= 12'd786;
            12'd54: PAGE <= 12'd1308;
            12'd55: PAGE <= 12'd1830;
            12'd56: PAGE <= 12'd299;
            12'd57: PAGE <= 12'd821;
            12'd58: PAGE <= 12'd1343;
            12'd59: PAGE <= 12'd1865;
            12'd60: PAGE <= 12'd334;
            12'd61: PAGE <= 12'd856;
            12'd62: PAGE <= 12'd1378;
            12'd63: PAGE <= 12'd1900;
            12'd64: PAGE <= 12'd369;
            12'd65: PAGE <= 12'd891;
            12'd66: PAGE <= 12'd1413;
            12'd67: PAGE <= 12'd1935;
            12'd68: PAGE <= 12'd404;
            12'd69: PAGE <= 12'd926;
            12'd70: PAGE <= 12'd1448;
            12'd71: PAGE <= 12'd1970;
            12'd72: PAGE <= 12'd439;
            12'd73: PAGE <= 12'd961;
            12'd74: PAGE <= 12'd1483;
            12'd75: PAGE <= 12'd2005;
            12'd76: PAGE <= 12'd474;
            12'd77: PAGE <= 12'd996;
            12'd78: PAGE <= 12'd1518;
            12'd79: PAGE <= 12'd2040;
            12'd80: PAGE <= 12'd509;
            12'd81: PAGE <= 12'd1031;
            12'd82: PAGE <= 12'd1553;
            12'd83: PAGE <= 12'd22;
            12'd84: PAGE <= 12'd544;
            12'd85: PAGE <= 12'd1066;
            12'd86: PAGE <= 12'd1588;
            12'd87: PAGE <= 12'd57;
            12'd88: PAGE <= 12'd579;
            12'd89: PAGE <= 12'd1101;
            12'd90: PAGE <= 12'd1623;
            12'd91: PAGE <= 12'd92;
            12'd92: PAGE <= 12'd614;
            12'd93: PAGE <= 12'd1136;
            12'd94: PAGE <= 12'd1658;
            12'd95: PAGE <= 12'd127;
            12'd96: PAGE <= 12'd649;
            12'd97: PAGE <= 12'd1171;
            12'd98: PAGE <= 12'd1693;
            12'd99: PAGE <= 12'd162;
            12'd100: PAGE <= 12'd684;
            12'd101: PAGE <= 12'd1206;
            12'd102: PAGE <= 12'd1728;
            12'd103: PAGE <= 12'd197;
            12'd104: PAGE <= 12'd719;
            12'd105: PAGE <= 12'd1241;
            12'd106: PAGE <= 12'd1763;
            12'd107: PAGE <= 12'd232;
            12'd108: PAGE <= 12'd754;
            12'd109: PAGE <= 12'd1276;
            12'd110: PAGE <= 12'd1798;
            12'd111: PAGE <= 12'd267;
            12'd112: PAGE <= 12'd789;
            12'd113: PAGE <= 12'd1311;
            12'd114: PAGE <= 12'd1833;
            12'd115: PAGE <= 12'd302;
            12'd116: PAGE <= 12'd824;
            12'd117: PAGE <= 12'd1346;
            12'd118: PAGE <= 12'd1868;
            12'd119: PAGE <= 12'd337;
            12'd120: PAGE <= 12'd859;
            12'd121: PAGE <= 12'd1381;
            12'd122: PAGE <= 12'd1903;
            12'd123: PAGE <= 12'd372;
            12'd124: PAGE <= 12'd894;
            12'd125: PAGE <= 12'd1416;
            12'd126: PAGE <= 12'd1938;
            12'd127: PAGE <= 12'd407;
            12'd128: PAGE <= 12'd929;
            12'd129: PAGE <= 12'd1451;
            12'd130: PAGE <= 12'd1973;
            12'd131: PAGE <= 12'd442;
            12'd132: PAGE <= 12'd964;
            12'd133: PAGE <= 12'd1486;
            12'd134: PAGE <= 12'd2008;
            12'd135: PAGE <= 12'd477;
            12'd136: PAGE <= 12'd999;
            12'd137: PAGE <= 12'd1521;
            12'd138: PAGE <= 12'd2043;
            12'd139: PAGE <= 12'd512;
            12'd140: PAGE <= 12'd1034;
            12'd141: PAGE <= 12'd1556;
            12'd142: PAGE <= 12'd25;
            12'd143: PAGE <= 12'd547;
            12'd144: PAGE <= 12'd1069;
            12'd145: PAGE <= 12'd1591;
            12'd146: PAGE <= 12'd60;
            12'd147: PAGE <= 12'd582;
            12'd148: PAGE <= 12'd1104;
            12'd149: PAGE <= 12'd1626;
            12'd150: PAGE <= 12'd95;
            12'd151: PAGE <= 12'd617;
            12'd152: PAGE <= 12'd1139;
            12'd153: PAGE <= 12'd1661;
            12'd154: PAGE <= 12'd130;
            12'd155: PAGE <= 12'd652;
            12'd156: PAGE <= 12'd1174;
            12'd157: PAGE <= 12'd1696;
            12'd158: PAGE <= 12'd165;
            12'd159: PAGE <= 12'd687;
            12'd160: PAGE <= 12'd1209;
            12'd161: PAGE <= 12'd1731;
            12'd162: PAGE <= 12'd200;
            12'd163: PAGE <= 12'd722;
            12'd164: PAGE <= 12'd1244;
            12'd165: PAGE <= 12'd1766;
            12'd166: PAGE <= 12'd235;
            12'd167: PAGE <= 12'd757;
            12'd168: PAGE <= 12'd1279;
            12'd169: PAGE <= 12'd1801;
            12'd170: PAGE <= 12'd270;
            12'd171: PAGE <= 12'd792;
            12'd172: PAGE <= 12'd1314;
            12'd173: PAGE <= 12'd1836;
            12'd174: PAGE <= 12'd305;
            12'd175: PAGE <= 12'd827;
            12'd176: PAGE <= 12'd1349;
            12'd177: PAGE <= 12'd1871;
            12'd178: PAGE <= 12'd340;
            12'd179: PAGE <= 12'd862;
            12'd180: PAGE <= 12'd1384;
            12'd181: PAGE <= 12'd1906;
            12'd182: PAGE <= 12'd375;
            12'd183: PAGE <= 12'd897;
            12'd184: PAGE <= 12'd1419;
            12'd185: PAGE <= 12'd1941;
            12'd186: PAGE <= 12'd410;
            12'd187: PAGE <= 12'd932;
            12'd188: PAGE <= 12'd1454;
            12'd189: PAGE <= 12'd1976;
            12'd190: PAGE <= 12'd445;
            12'd191: PAGE <= 12'd967;
            12'd192: PAGE <= 12'd1489;
            12'd193: PAGE <= 12'd2011;
            12'd194: PAGE <= 12'd480;
            12'd195: PAGE <= 12'd1002;
            12'd196: PAGE <= 12'd1524;
            12'd197: PAGE <= 12'd2046;
            12'd198: PAGE <= 12'd515;
            12'd199: PAGE <= 12'd1037;
            12'd200: PAGE <= 12'd1559;
            12'd201: PAGE <= 12'd28;
            12'd202: PAGE <= 12'd550;
            12'd203: PAGE <= 12'd1072;
            12'd204: PAGE <= 12'd1594;
            12'd205: PAGE <= 12'd63;
            12'd206: PAGE <= 12'd585;
            12'd207: PAGE <= 12'd1107;
            12'd208: PAGE <= 12'd1629;
            12'd209: PAGE <= 12'd98;
            12'd210: PAGE <= 12'd620;
            12'd211: PAGE <= 12'd1142;
            12'd212: PAGE <= 12'd1664;
            12'd213: PAGE <= 12'd133;
            12'd214: PAGE <= 12'd655;
            12'd215: PAGE <= 12'd1177;
            12'd216: PAGE <= 12'd1699;
            12'd217: PAGE <= 12'd168;
            12'd218: PAGE <= 12'd690;
            12'd219: PAGE <= 12'd1212;
            12'd220: PAGE <= 12'd1734;
            12'd221: PAGE <= 12'd203;
            12'd222: PAGE <= 12'd725;
            12'd223: PAGE <= 12'd1247;
            12'd224: PAGE <= 12'd1769;
            12'd225: PAGE <= 12'd238;
            12'd226: PAGE <= 12'd760;
            12'd227: PAGE <= 12'd1282;
            12'd228: PAGE <= 12'd1804;
            12'd229: PAGE <= 12'd273;
            12'd230: PAGE <= 12'd795;
            12'd231: PAGE <= 12'd1317;
            12'd232: PAGE <= 12'd1839;
            12'd233: PAGE <= 12'd308;
            12'd234: PAGE <= 12'd830;
            12'd235: PAGE <= 12'd1352;
            12'd236: PAGE <= 12'd1874;
            12'd237: PAGE <= 12'd343;
            12'd238: PAGE <= 12'd865;
            12'd239: PAGE <= 12'd1387;
            12'd240: PAGE <= 12'd1909;
            12'd241: PAGE <= 12'd378;
            12'd242: PAGE <= 12'd900;
            12'd243: PAGE <= 12'd1422;
            12'd244: PAGE <= 12'd1944;
            12'd245: PAGE <= 12'd413;
            12'd246: PAGE <= 12'd935;
            12'd247: PAGE <= 12'd1457;
            12'd248: PAGE <= 12'd1979;
            12'd249: PAGE <= 12'd448;
            12'd250: PAGE <= 12'd970;
            12'd251: PAGE <= 12'd1492;
            12'd252: PAGE <= 12'd2014;
            12'd253: PAGE <= 12'd483;
            12'd254: PAGE <= 12'd1005;
            12'd255: PAGE <= 12'd1527;
            12'd256: PAGE <= 12'd2049;
            12'd257: PAGE <= 12'd518;
            12'd258: PAGE <= 12'd1040;
            12'd259: PAGE <= 12'd1562;
            12'd260: PAGE <= 12'd31;
            12'd261: PAGE <= 12'd553;
            12'd262: PAGE <= 12'd1075;
            12'd263: PAGE <= 12'd1597;
            12'd264: PAGE <= 12'd66;
            12'd265: PAGE <= 12'd588;
            12'd266: PAGE <= 12'd1110;
            12'd267: PAGE <= 12'd1632;
            12'd268: PAGE <= 12'd101;
            12'd269: PAGE <= 12'd623;
            12'd270: PAGE <= 12'd1145;
            12'd271: PAGE <= 12'd1667;
            12'd272: PAGE <= 12'd136;
            12'd273: PAGE <= 12'd658;
            12'd274: PAGE <= 12'd1180;
            12'd275: PAGE <= 12'd1702;
            12'd276: PAGE <= 12'd171;
            12'd277: PAGE <= 12'd693;
            12'd278: PAGE <= 12'd1215;
            12'd279: PAGE <= 12'd1737;
            12'd280: PAGE <= 12'd206;
            12'd281: PAGE <= 12'd728;
            12'd282: PAGE <= 12'd1250;
            12'd283: PAGE <= 12'd1772;
            12'd284: PAGE <= 12'd241;
            12'd285: PAGE <= 12'd763;
            12'd286: PAGE <= 12'd1285;
            12'd287: PAGE <= 12'd1807;
            12'd288: PAGE <= 12'd276;
            12'd289: PAGE <= 12'd798;
            12'd290: PAGE <= 12'd1320;
            12'd291: PAGE <= 12'd1842;
            12'd292: PAGE <= 12'd311;
            12'd293: PAGE <= 12'd833;
            12'd294: PAGE <= 12'd1355;
            12'd295: PAGE <= 12'd1877;
            12'd296: PAGE <= 12'd346;
            12'd297: PAGE <= 12'd868;
            12'd298: PAGE <= 12'd1390;
            12'd299: PAGE <= 12'd1912;
            12'd300: PAGE <= 12'd381;
            12'd301: PAGE <= 12'd903;
            12'd302: PAGE <= 12'd1425;
            12'd303: PAGE <= 12'd1947;
            12'd304: PAGE <= 12'd416;
            12'd305: PAGE <= 12'd938;
            12'd306: PAGE <= 12'd1460;
            12'd307: PAGE <= 12'd1982;
            12'd308: PAGE <= 12'd451;
            12'd309: PAGE <= 12'd973;
            12'd310: PAGE <= 12'd1495;
            12'd311: PAGE <= 12'd2017;
            12'd312: PAGE <= 12'd486;
            12'd313: PAGE <= 12'd1008;
            12'd314: PAGE <= 12'd1530;
            12'd315: PAGE <= 12'd2052;
            12'd316: PAGE <= 12'd521;
            12'd317: PAGE <= 12'd1043;
            12'd318: PAGE <= 12'd1565;
            12'd319: PAGE <= 12'd34;
            12'd320: PAGE <= 12'd556;
            12'd321: PAGE <= 12'd1078;
            12'd322: PAGE <= 12'd1600;
            12'd323: PAGE <= 12'd69;
            12'd324: PAGE <= 12'd591;
            12'd325: PAGE <= 12'd1113;
            12'd326: PAGE <= 12'd1635;
            12'd327: PAGE <= 12'd104;
            12'd328: PAGE <= 12'd626;
            12'd329: PAGE <= 12'd1148;
            12'd330: PAGE <= 12'd1670;
            12'd331: PAGE <= 12'd139;
            12'd332: PAGE <= 12'd661;
            12'd333: PAGE <= 12'd1183;
            12'd334: PAGE <= 12'd1705;
            12'd335: PAGE <= 12'd174;
            12'd336: PAGE <= 12'd696;
            12'd337: PAGE <= 12'd1218;
            12'd338: PAGE <= 12'd1740;
            12'd339: PAGE <= 12'd209;
            12'd340: PAGE <= 12'd731;
            12'd341: PAGE <= 12'd1253;
            12'd342: PAGE <= 12'd1775;
            12'd343: PAGE <= 12'd244;
            12'd344: PAGE <= 12'd766;
            12'd345: PAGE <= 12'd1288;
            12'd346: PAGE <= 12'd1810;
            12'd347: PAGE <= 12'd279;
            12'd348: PAGE <= 12'd801;
            12'd349: PAGE <= 12'd1323;
            12'd350: PAGE <= 12'd1845;
            12'd351: PAGE <= 12'd314;
            12'd352: PAGE <= 12'd836;
            12'd353: PAGE <= 12'd1358;
            12'd354: PAGE <= 12'd1880;
            12'd355: PAGE <= 12'd349;
            12'd356: PAGE <= 12'd871;
            12'd357: PAGE <= 12'd1393;
            12'd358: PAGE <= 12'd1915;
            12'd359: PAGE <= 12'd384;
            12'd360: PAGE <= 12'd906;
            12'd361: PAGE <= 12'd1428;
            12'd362: PAGE <= 12'd1950;
            12'd363: PAGE <= 12'd419;
            12'd364: PAGE <= 12'd941;
            12'd365: PAGE <= 12'd1463;
            12'd366: PAGE <= 12'd1985;
            12'd367: PAGE <= 12'd454;
            12'd368: PAGE <= 12'd976;
            12'd369: PAGE <= 12'd1498;
            12'd370: PAGE <= 12'd2020;
            12'd371: PAGE <= 12'd489;
            12'd372: PAGE <= 12'd1011;
            12'd373: PAGE <= 12'd1533;
            12'd374: PAGE <= 12'd2;
            12'd375: PAGE <= 12'd524;
            12'd376: PAGE <= 12'd1046;
            12'd377: PAGE <= 12'd1568;
            12'd378: PAGE <= 12'd37;
            12'd379: PAGE <= 12'd559;
            12'd380: PAGE <= 12'd1081;
            12'd381: PAGE <= 12'd1603;
            12'd382: PAGE <= 12'd72;
            12'd383: PAGE <= 12'd594;
            12'd384: PAGE <= 12'd1116;
            12'd385: PAGE <= 12'd1638;
            12'd386: PAGE <= 12'd107;
            12'd387: PAGE <= 12'd629;
            12'd388: PAGE <= 12'd1151;
            12'd389: PAGE <= 12'd1673;
            12'd390: PAGE <= 12'd142;
            12'd391: PAGE <= 12'd664;
            12'd392: PAGE <= 12'd1186;
            12'd393: PAGE <= 12'd1708;
            12'd394: PAGE <= 12'd177;
            12'd395: PAGE <= 12'd699;
            12'd396: PAGE <= 12'd1221;
            12'd397: PAGE <= 12'd1743;
            12'd398: PAGE <= 12'd212;
            12'd399: PAGE <= 12'd734;
            12'd400: PAGE <= 12'd1256;
            12'd401: PAGE <= 12'd1778;
            12'd402: PAGE <= 12'd247;
            12'd403: PAGE <= 12'd769;
            12'd404: PAGE <= 12'd1291;
            12'd405: PAGE <= 12'd1813;
            12'd406: PAGE <= 12'd282;
            12'd407: PAGE <= 12'd804;
            12'd408: PAGE <= 12'd1326;
            12'd409: PAGE <= 12'd1848;
            12'd410: PAGE <= 12'd317;
            12'd411: PAGE <= 12'd839;
            12'd412: PAGE <= 12'd1361;
            12'd413: PAGE <= 12'd1883;
            12'd414: PAGE <= 12'd352;
            12'd415: PAGE <= 12'd874;
            12'd416: PAGE <= 12'd1396;
            12'd417: PAGE <= 12'd1918;
            12'd418: PAGE <= 12'd387;
            12'd419: PAGE <= 12'd909;
            12'd420: PAGE <= 12'd1431;
            12'd421: PAGE <= 12'd1953;
            12'd422: PAGE <= 12'd422;
            12'd423: PAGE <= 12'd944;
            12'd424: PAGE <= 12'd1466;
            12'd425: PAGE <= 12'd1988;
            12'd426: PAGE <= 12'd457;
            12'd427: PAGE <= 12'd979;
            12'd428: PAGE <= 12'd1501;
            12'd429: PAGE <= 12'd2023;
            12'd430: PAGE <= 12'd492;
            12'd431: PAGE <= 12'd1014;
            12'd432: PAGE <= 12'd1536;
            12'd433: PAGE <= 12'd5;
            12'd434: PAGE <= 12'd527;
            12'd435: PAGE <= 12'd1049;
            12'd436: PAGE <= 12'd1571;
            12'd437: PAGE <= 12'd40;
            12'd438: PAGE <= 12'd562;
            12'd439: PAGE <= 12'd1084;
            12'd440: PAGE <= 12'd1606;
            12'd441: PAGE <= 12'd75;
            12'd442: PAGE <= 12'd597;
            12'd443: PAGE <= 12'd1119;
            12'd444: PAGE <= 12'd1641;
            12'd445: PAGE <= 12'd110;
            12'd446: PAGE <= 12'd632;
            12'd447: PAGE <= 12'd1154;
            12'd448: PAGE <= 12'd1676;
            12'd449: PAGE <= 12'd145;
            12'd450: PAGE <= 12'd667;
            12'd451: PAGE <= 12'd1189;
            12'd452: PAGE <= 12'd1711;
            12'd453: PAGE <= 12'd180;
            12'd454: PAGE <= 12'd702;
            12'd455: PAGE <= 12'd1224;
            12'd456: PAGE <= 12'd1746;
            12'd457: PAGE <= 12'd215;
            12'd458: PAGE <= 12'd737;
            12'd459: PAGE <= 12'd1259;
            12'd460: PAGE <= 12'd1781;
            12'd461: PAGE <= 12'd250;
            12'd462: PAGE <= 12'd772;
            12'd463: PAGE <= 12'd1294;
            12'd464: PAGE <= 12'd1816;
            12'd465: PAGE <= 12'd285;
            12'd466: PAGE <= 12'd807;
            12'd467: PAGE <= 12'd1329;
            12'd468: PAGE <= 12'd1851;
            12'd469: PAGE <= 12'd320;
            12'd470: PAGE <= 12'd842;
            12'd471: PAGE <= 12'd1364;
            12'd472: PAGE <= 12'd1886;
            12'd473: PAGE <= 12'd355;
            12'd474: PAGE <= 12'd877;
            12'd475: PAGE <= 12'd1399;
            12'd476: PAGE <= 12'd1921;
            12'd477: PAGE <= 12'd390;
            12'd478: PAGE <= 12'd912;
            12'd479: PAGE <= 12'd1434;
            12'd480: PAGE <= 12'd1956;
            12'd481: PAGE <= 12'd425;
            12'd482: PAGE <= 12'd947;
            12'd483: PAGE <= 12'd1469;
            12'd484: PAGE <= 12'd1991;
            12'd485: PAGE <= 12'd460;
            12'd486: PAGE <= 12'd982;
            12'd487: PAGE <= 12'd1504;
            12'd488: PAGE <= 12'd2026;
            12'd489: PAGE <= 12'd495;
            12'd490: PAGE <= 12'd1017;
            12'd491: PAGE <= 12'd1539;
            12'd492: PAGE <= 12'd8;
            12'd493: PAGE <= 12'd530;
            12'd494: PAGE <= 12'd1052;
            12'd495: PAGE <= 12'd1574;
            12'd496: PAGE <= 12'd43;
            12'd497: PAGE <= 12'd565;
            12'd498: PAGE <= 12'd1087;
            12'd499: PAGE <= 12'd1609;
            12'd500: PAGE <= 12'd78;
            12'd501: PAGE <= 12'd600;
            12'd502: PAGE <= 12'd1122;
            12'd503: PAGE <= 12'd1644;
            12'd504: PAGE <= 12'd113;
            12'd505: PAGE <= 12'd635;
            12'd506: PAGE <= 12'd1157;
            12'd507: PAGE <= 12'd1679;
            12'd508: PAGE <= 12'd148;
            12'd509: PAGE <= 12'd670;
            12'd510: PAGE <= 12'd1192;
            12'd511: PAGE <= 12'd1714;
            12'd512: PAGE <= 12'd183;
            12'd513: PAGE <= 12'd705;
            12'd514: PAGE <= 12'd1227;
            12'd515: PAGE <= 12'd1749;
            12'd516: PAGE <= 12'd218;
            12'd517: PAGE <= 12'd740;
            12'd518: PAGE <= 12'd1262;
            12'd519: PAGE <= 12'd1784;
            12'd520: PAGE <= 12'd253;
            12'd521: PAGE <= 12'd775;
            12'd522: PAGE <= 12'd1297;
            12'd523: PAGE <= 12'd1819;
            12'd524: PAGE <= 12'd288;
            12'd525: PAGE <= 12'd810;
            12'd526: PAGE <= 12'd1332;
            12'd527: PAGE <= 12'd1854;
            12'd528: PAGE <= 12'd323;
            12'd529: PAGE <= 12'd845;
            12'd530: PAGE <= 12'd1367;
            12'd531: PAGE <= 12'd1889;
            12'd532: PAGE <= 12'd358;
            12'd533: PAGE <= 12'd880;
            12'd534: PAGE <= 12'd1402;
            12'd535: PAGE <= 12'd1924;
            12'd536: PAGE <= 12'd393;
            12'd537: PAGE <= 12'd915;
            12'd538: PAGE <= 12'd1437;
            12'd539: PAGE <= 12'd1959;
            12'd540: PAGE <= 12'd428;
            12'd541: PAGE <= 12'd950;
            12'd542: PAGE <= 12'd1472;
            12'd543: PAGE <= 12'd1994;
            12'd544: PAGE <= 12'd463;
            12'd545: PAGE <= 12'd985;
            12'd546: PAGE <= 12'd1507;
            12'd547: PAGE <= 12'd2029;
            12'd548: PAGE <= 12'd498;
            12'd549: PAGE <= 12'd1020;
            12'd550: PAGE <= 12'd1542;
            12'd551: PAGE <= 12'd11;
            12'd552: PAGE <= 12'd533;
            12'd553: PAGE <= 12'd1055;
            12'd554: PAGE <= 12'd1577;
            12'd555: PAGE <= 12'd46;
            12'd556: PAGE <= 12'd568;
            12'd557: PAGE <= 12'd1090;
            12'd558: PAGE <= 12'd1612;
            12'd559: PAGE <= 12'd81;
            12'd560: PAGE <= 12'd603;
            12'd561: PAGE <= 12'd1125;
            12'd562: PAGE <= 12'd1647;
            12'd563: PAGE <= 12'd116;
            12'd564: PAGE <= 12'd638;
            12'd565: PAGE <= 12'd1160;
            12'd566: PAGE <= 12'd1682;
            12'd567: PAGE <= 12'd151;
            12'd568: PAGE <= 12'd673;
            12'd569: PAGE <= 12'd1195;
            12'd570: PAGE <= 12'd1717;
            12'd571: PAGE <= 12'd186;
            12'd572: PAGE <= 12'd708;
            12'd573: PAGE <= 12'd1230;
            12'd574: PAGE <= 12'd1752;
            12'd575: PAGE <= 12'd221;
            12'd576: PAGE <= 12'd743;
            12'd577: PAGE <= 12'd1265;
            12'd578: PAGE <= 12'd1787;
            12'd579: PAGE <= 12'd256;
            12'd580: PAGE <= 12'd778;
            12'd581: PAGE <= 12'd1300;
            12'd582: PAGE <= 12'd1822;
            12'd583: PAGE <= 12'd291;
            12'd584: PAGE <= 12'd813;
            12'd585: PAGE <= 12'd1335;
            12'd586: PAGE <= 12'd1857;
            12'd587: PAGE <= 12'd326;
            12'd588: PAGE <= 12'd848;
            12'd589: PAGE <= 12'd1370;
            12'd590: PAGE <= 12'd1892;
            12'd591: PAGE <= 12'd361;
            12'd592: PAGE <= 12'd883;
            12'd593: PAGE <= 12'd1405;
            12'd594: PAGE <= 12'd1927;
            12'd595: PAGE <= 12'd396;
            12'd596: PAGE <= 12'd918;
            12'd597: PAGE <= 12'd1440;
            12'd598: PAGE <= 12'd1962;
            12'd599: PAGE <= 12'd431;
            12'd600: PAGE <= 12'd953;
            12'd601: PAGE <= 12'd1475;
            12'd602: PAGE <= 12'd1997;
            12'd603: PAGE <= 12'd466;
            12'd604: PAGE <= 12'd988;
            12'd605: PAGE <= 12'd1510;
            12'd606: PAGE <= 12'd2032;
            12'd607: PAGE <= 12'd501;
            12'd608: PAGE <= 12'd1023;
            12'd609: PAGE <= 12'd1545;
            12'd610: PAGE <= 12'd14;
            12'd611: PAGE <= 12'd536;
            12'd612: PAGE <= 12'd1058;
            12'd613: PAGE <= 12'd1580;
            12'd614: PAGE <= 12'd49;
            12'd615: PAGE <= 12'd571;
            12'd616: PAGE <= 12'd1093;
            12'd617: PAGE <= 12'd1615;
            12'd618: PAGE <= 12'd84;
            12'd619: PAGE <= 12'd606;
            12'd620: PAGE <= 12'd1128;
            12'd621: PAGE <= 12'd1650;
            12'd622: PAGE <= 12'd119;
            12'd623: PAGE <= 12'd641;
            12'd624: PAGE <= 12'd1163;
            12'd625: PAGE <= 12'd1685;
            12'd626: PAGE <= 12'd154;
            12'd627: PAGE <= 12'd676;
            12'd628: PAGE <= 12'd1198;
            12'd629: PAGE <= 12'd1720;
            12'd630: PAGE <= 12'd189;
            12'd631: PAGE <= 12'd711;
            12'd632: PAGE <= 12'd1233;
            12'd633: PAGE <= 12'd1755;
            12'd634: PAGE <= 12'd224;
            12'd635: PAGE <= 12'd746;
            12'd636: PAGE <= 12'd1268;
            12'd637: PAGE <= 12'd1790;
            12'd638: PAGE <= 12'd259;
            12'd639: PAGE <= 12'd781;
            12'd640: PAGE <= 12'd1303;
            12'd641: PAGE <= 12'd1825;
            12'd642: PAGE <= 12'd294;
            12'd643: PAGE <= 12'd816;
            12'd644: PAGE <= 12'd1338;
            12'd645: PAGE <= 12'd1860;
            12'd646: PAGE <= 12'd329;
            12'd647: PAGE <= 12'd851;
            12'd648: PAGE <= 12'd1373;
            12'd649: PAGE <= 12'd1895;
            12'd650: PAGE <= 12'd364;
            12'd651: PAGE <= 12'd886;
            12'd652: PAGE <= 12'd1408;
            12'd653: PAGE <= 12'd1930;
            12'd654: PAGE <= 12'd399;
            12'd655: PAGE <= 12'd921;
            12'd656: PAGE <= 12'd1443;
            12'd657: PAGE <= 12'd1965;
            12'd658: PAGE <= 12'd434;
            12'd659: PAGE <= 12'd956;
            12'd660: PAGE <= 12'd1478;
            12'd661: PAGE <= 12'd2000;
            12'd662: PAGE <= 12'd469;
            12'd663: PAGE <= 12'd991;
            12'd664: PAGE <= 12'd1513;
            12'd665: PAGE <= 12'd2035;
            12'd666: PAGE <= 12'd504;
            12'd667: PAGE <= 12'd1026;
            12'd668: PAGE <= 12'd1548;
            12'd669: PAGE <= 12'd17;
            12'd670: PAGE <= 12'd539;
            12'd671: PAGE <= 12'd1061;
            12'd672: PAGE <= 12'd1583;
            12'd673: PAGE <= 12'd52;
            12'd674: PAGE <= 12'd574;
            12'd675: PAGE <= 12'd1096;
            12'd676: PAGE <= 12'd1618;
            12'd677: PAGE <= 12'd87;
            12'd678: PAGE <= 12'd609;
            12'd679: PAGE <= 12'd1131;
            12'd680: PAGE <= 12'd1653;
            12'd681: PAGE <= 12'd122;
            12'd682: PAGE <= 12'd644;
            12'd683: PAGE <= 12'd1166;
            12'd684: PAGE <= 12'd1688;
            12'd685: PAGE <= 12'd157;
            12'd686: PAGE <= 12'd679;
            12'd687: PAGE <= 12'd1201;
            12'd688: PAGE <= 12'd1723;
            12'd689: PAGE <= 12'd192;
            12'd690: PAGE <= 12'd714;
            12'd691: PAGE <= 12'd1236;
            12'd692: PAGE <= 12'd1758;
            12'd693: PAGE <= 12'd227;
            12'd694: PAGE <= 12'd749;
            12'd695: PAGE <= 12'd1271;
            12'd696: PAGE <= 12'd1793;
            12'd697: PAGE <= 12'd262;
            12'd698: PAGE <= 12'd784;
            12'd699: PAGE <= 12'd1306;
            12'd700: PAGE <= 12'd1828;
            12'd701: PAGE <= 12'd297;
            12'd702: PAGE <= 12'd819;
            12'd703: PAGE <= 12'd1341;
            12'd704: PAGE <= 12'd1863;
            12'd705: PAGE <= 12'd332;
            12'd706: PAGE <= 12'd854;
            12'd707: PAGE <= 12'd1376;
            12'd708: PAGE <= 12'd1898;
            12'd709: PAGE <= 12'd367;
            12'd710: PAGE <= 12'd889;
            12'd711: PAGE <= 12'd1411;
            12'd712: PAGE <= 12'd1933;
            12'd713: PAGE <= 12'd402;
            12'd714: PAGE <= 12'd924;
            12'd715: PAGE <= 12'd1446;
            12'd716: PAGE <= 12'd1968;
            12'd717: PAGE <= 12'd437;
            12'd718: PAGE <= 12'd959;
            12'd719: PAGE <= 12'd1481;
            12'd720: PAGE <= 12'd2003;
            12'd721: PAGE <= 12'd472;
            12'd722: PAGE <= 12'd994;
            12'd723: PAGE <= 12'd1516;
            12'd724: PAGE <= 12'd2038;
            12'd725: PAGE <= 12'd507;
            12'd726: PAGE <= 12'd1029;
            12'd727: PAGE <= 12'd1551;
            12'd728: PAGE <= 12'd20;
            12'd729: PAGE <= 12'd542;
            12'd730: PAGE <= 12'd1064;
            12'd731: PAGE <= 12'd1586;
            12'd732: PAGE <= 12'd55;
            12'd733: PAGE <= 12'd577;
            12'd734: PAGE <= 12'd1099;
            12'd735: PAGE <= 12'd1621;
            12'd736: PAGE <= 12'd90;
            12'd737: PAGE <= 12'd612;
            12'd738: PAGE <= 12'd1134;
            12'd739: PAGE <= 12'd1656;
            12'd740: PAGE <= 12'd125;
            12'd741: PAGE <= 12'd647;
            12'd742: PAGE <= 12'd1169;
            12'd743: PAGE <= 12'd1691;
            12'd744: PAGE <= 12'd160;
            12'd745: PAGE <= 12'd682;
            12'd746: PAGE <= 12'd1204;
            12'd747: PAGE <= 12'd1726;
            12'd748: PAGE <= 12'd195;
            12'd749: PAGE <= 12'd717;
            12'd750: PAGE <= 12'd1239;
            12'd751: PAGE <= 12'd1761;
            12'd752: PAGE <= 12'd230;
            12'd753: PAGE <= 12'd752;
            12'd754: PAGE <= 12'd1274;
            12'd755: PAGE <= 12'd1796;
            12'd756: PAGE <= 12'd265;
            12'd757: PAGE <= 12'd787;
            12'd758: PAGE <= 12'd1309;
            12'd759: PAGE <= 12'd1831;
            12'd760: PAGE <= 12'd300;
            12'd761: PAGE <= 12'd822;
            12'd762: PAGE <= 12'd1344;
            12'd763: PAGE <= 12'd1866;
            12'd764: PAGE <= 12'd335;
            12'd765: PAGE <= 12'd857;
            12'd766: PAGE <= 12'd1379;
            12'd767: PAGE <= 12'd1901;
            12'd768: PAGE <= 12'd370;
            12'd769: PAGE <= 12'd892;
            12'd770: PAGE <= 12'd1414;
            12'd771: PAGE <= 12'd1936;
            12'd772: PAGE <= 12'd405;
            12'd773: PAGE <= 12'd927;
            12'd774: PAGE <= 12'd1449;
            12'd775: PAGE <= 12'd1971;
            12'd776: PAGE <= 12'd440;
            12'd777: PAGE <= 12'd962;
            12'd778: PAGE <= 12'd1484;
            12'd779: PAGE <= 12'd2006;
            12'd780: PAGE <= 12'd475;
            12'd781: PAGE <= 12'd997;
            12'd782: PAGE <= 12'd1519;
            12'd783: PAGE <= 12'd2041;
            12'd784: PAGE <= 12'd510;
            12'd785: PAGE <= 12'd1032;
            12'd786: PAGE <= 12'd1554;
            12'd787: PAGE <= 12'd23;
            12'd788: PAGE <= 12'd545;
            12'd789: PAGE <= 12'd1067;
            12'd790: PAGE <= 12'd1589;
            12'd791: PAGE <= 12'd58;
            12'd792: PAGE <= 12'd580;
            12'd793: PAGE <= 12'd1102;
            12'd794: PAGE <= 12'd1624;
            12'd795: PAGE <= 12'd93;
            12'd796: PAGE <= 12'd615;
            12'd797: PAGE <= 12'd1137;
            12'd798: PAGE <= 12'd1659;
            12'd799: PAGE <= 12'd128;
            12'd800: PAGE <= 12'd650;
            12'd801: PAGE <= 12'd1172;
            12'd802: PAGE <= 12'd1694;
            12'd803: PAGE <= 12'd163;
            12'd804: PAGE <= 12'd685;
            12'd805: PAGE <= 12'd1207;
            12'd806: PAGE <= 12'd1729;
            12'd807: PAGE <= 12'd198;
            12'd808: PAGE <= 12'd720;
            12'd809: PAGE <= 12'd1242;
            12'd810: PAGE <= 12'd1764;
            12'd811: PAGE <= 12'd233;
            12'd812: PAGE <= 12'd755;
            12'd813: PAGE <= 12'd1277;
            12'd814: PAGE <= 12'd1799;
            12'd815: PAGE <= 12'd268;
            12'd816: PAGE <= 12'd790;
            12'd817: PAGE <= 12'd1312;
            12'd818: PAGE <= 12'd1834;
            12'd819: PAGE <= 12'd303;
            12'd820: PAGE <= 12'd825;
            12'd821: PAGE <= 12'd1347;
            12'd822: PAGE <= 12'd1869;
            12'd823: PAGE <= 12'd338;
            12'd824: PAGE <= 12'd860;
            12'd825: PAGE <= 12'd1382;
            12'd826: PAGE <= 12'd1904;
            12'd827: PAGE <= 12'd373;
            12'd828: PAGE <= 12'd895;
            12'd829: PAGE <= 12'd1417;
            12'd830: PAGE <= 12'd1939;
            12'd831: PAGE <= 12'd408;
            12'd832: PAGE <= 12'd930;
            12'd833: PAGE <= 12'd1452;
            12'd834: PAGE <= 12'd1974;
            12'd835: PAGE <= 12'd443;
            12'd836: PAGE <= 12'd965;
            12'd837: PAGE <= 12'd1487;
            12'd838: PAGE <= 12'd2009;
            12'd839: PAGE <= 12'd478;
            12'd840: PAGE <= 12'd1000;
            12'd841: PAGE <= 12'd1522;
            12'd842: PAGE <= 12'd2044;
            12'd843: PAGE <= 12'd513;
            12'd844: PAGE <= 12'd1035;
            12'd845: PAGE <= 12'd1557;
            12'd846: PAGE <= 12'd26;
            12'd847: PAGE <= 12'd548;
            12'd848: PAGE <= 12'd1070;
            12'd849: PAGE <= 12'd1592;
            12'd850: PAGE <= 12'd61;
            12'd851: PAGE <= 12'd583;
            12'd852: PAGE <= 12'd1105;
            12'd853: PAGE <= 12'd1627;
            12'd854: PAGE <= 12'd96;
            12'd855: PAGE <= 12'd618;
            12'd856: PAGE <= 12'd1140;
            12'd857: PAGE <= 12'd1662;
            12'd858: PAGE <= 12'd131;
            12'd859: PAGE <= 12'd653;
            12'd860: PAGE <= 12'd1175;
            12'd861: PAGE <= 12'd1697;
            12'd862: PAGE <= 12'd166;
            12'd863: PAGE <= 12'd688;
            12'd864: PAGE <= 12'd1210;
            12'd865: PAGE <= 12'd1732;
            12'd866: PAGE <= 12'd201;
            12'd867: PAGE <= 12'd723;
            12'd868: PAGE <= 12'd1245;
            12'd869: PAGE <= 12'd1767;
            12'd870: PAGE <= 12'd236;
            12'd871: PAGE <= 12'd758;
            12'd872: PAGE <= 12'd1280;
            12'd873: PAGE <= 12'd1802;
            12'd874: PAGE <= 12'd271;
            12'd875: PAGE <= 12'd793;
            12'd876: PAGE <= 12'd1315;
            12'd877: PAGE <= 12'd1837;
            12'd878: PAGE <= 12'd306;
            12'd879: PAGE <= 12'd828;
            12'd880: PAGE <= 12'd1350;
            12'd881: PAGE <= 12'd1872;
            12'd882: PAGE <= 12'd341;
            12'd883: PAGE <= 12'd863;
            12'd884: PAGE <= 12'd1385;
            12'd885: PAGE <= 12'd1907;
            12'd886: PAGE <= 12'd376;
            12'd887: PAGE <= 12'd898;
            12'd888: PAGE <= 12'd1420;
            12'd889: PAGE <= 12'd1942;
            12'd890: PAGE <= 12'd411;
            12'd891: PAGE <= 12'd933;
            12'd892: PAGE <= 12'd1455;
            12'd893: PAGE <= 12'd1977;
            12'd894: PAGE <= 12'd446;
            12'd895: PAGE <= 12'd968;
            12'd896: PAGE <= 12'd1490;
            12'd897: PAGE <= 12'd2012;
            12'd898: PAGE <= 12'd481;
            12'd899: PAGE <= 12'd1003;
            12'd900: PAGE <= 12'd1525;
            12'd901: PAGE <= 12'd2047;
            12'd902: PAGE <= 12'd516;
            12'd903: PAGE <= 12'd1038;
            12'd904: PAGE <= 12'd1560;
            12'd905: PAGE <= 12'd29;
            12'd906: PAGE <= 12'd551;
            12'd907: PAGE <= 12'd1073;
            12'd908: PAGE <= 12'd1595;
            12'd909: PAGE <= 12'd64;
            12'd910: PAGE <= 12'd586;
            12'd911: PAGE <= 12'd1108;
            12'd912: PAGE <= 12'd1630;
            12'd913: PAGE <= 12'd99;
            12'd914: PAGE <= 12'd621;
            12'd915: PAGE <= 12'd1143;
            12'd916: PAGE <= 12'd1665;
            12'd917: PAGE <= 12'd134;
            12'd918: PAGE <= 12'd656;
            12'd919: PAGE <= 12'd1178;
            12'd920: PAGE <= 12'd1700;
            12'd921: PAGE <= 12'd169;
            12'd922: PAGE <= 12'd691;
            12'd923: PAGE <= 12'd1213;
            12'd924: PAGE <= 12'd1735;
            12'd925: PAGE <= 12'd204;
            12'd926: PAGE <= 12'd726;
            12'd927: PAGE <= 12'd1248;
            12'd928: PAGE <= 12'd1770;
            12'd929: PAGE <= 12'd239;
            12'd930: PAGE <= 12'd761;
            12'd931: PAGE <= 12'd1283;
            12'd932: PAGE <= 12'd1805;
            12'd933: PAGE <= 12'd274;
            12'd934: PAGE <= 12'd796;
            12'd935: PAGE <= 12'd1318;
            12'd936: PAGE <= 12'd1840;
            12'd937: PAGE <= 12'd309;
            12'd938: PAGE <= 12'd831;
            12'd939: PAGE <= 12'd1353;
            12'd940: PAGE <= 12'd1875;
            12'd941: PAGE <= 12'd344;
            12'd942: PAGE <= 12'd866;
            12'd943: PAGE <= 12'd1388;
            12'd944: PAGE <= 12'd1910;
            12'd945: PAGE <= 12'd379;
            12'd946: PAGE <= 12'd901;
            12'd947: PAGE <= 12'd1423;
            12'd948: PAGE <= 12'd1945;
            12'd949: PAGE <= 12'd414;
            12'd950: PAGE <= 12'd936;
            12'd951: PAGE <= 12'd1458;
            12'd952: PAGE <= 12'd1980;
            12'd953: PAGE <= 12'd449;
            12'd954: PAGE <= 12'd971;
            12'd955: PAGE <= 12'd1493;
            12'd956: PAGE <= 12'd2015;
            12'd957: PAGE <= 12'd484;
            12'd958: PAGE <= 12'd1006;
            12'd959: PAGE <= 12'd1528;
            12'd960: PAGE <= 12'd2050;
            12'd961: PAGE <= 12'd519;
            12'd962: PAGE <= 12'd1041;
            12'd963: PAGE <= 12'd1563;
            12'd964: PAGE <= 12'd32;
            12'd965: PAGE <= 12'd554;
            12'd966: PAGE <= 12'd1076;
            12'd967: PAGE <= 12'd1598;
            12'd968: PAGE <= 12'd67;
            12'd969: PAGE <= 12'd589;
            12'd970: PAGE <= 12'd1111;
            12'd971: PAGE <= 12'd1633;
            12'd972: PAGE <= 12'd102;
            12'd973: PAGE <= 12'd624;
            12'd974: PAGE <= 12'd1146;
            12'd975: PAGE <= 12'd1668;
            12'd976: PAGE <= 12'd137;
            12'd977: PAGE <= 12'd659;
            12'd978: PAGE <= 12'd1181;
            12'd979: PAGE <= 12'd1703;
            12'd980: PAGE <= 12'd172;
            12'd981: PAGE <= 12'd694;
            12'd982: PAGE <= 12'd1216;
            12'd983: PAGE <= 12'd1738;
            12'd984: PAGE <= 12'd207;
            12'd985: PAGE <= 12'd729;
            12'd986: PAGE <= 12'd1251;
            12'd987: PAGE <= 12'd1773;
            12'd988: PAGE <= 12'd242;
            12'd989: PAGE <= 12'd764;
            12'd990: PAGE <= 12'd1286;
            12'd991: PAGE <= 12'd1808;
            12'd992: PAGE <= 12'd277;
            12'd993: PAGE <= 12'd799;
            12'd994: PAGE <= 12'd1321;
            12'd995: PAGE <= 12'd1843;
            12'd996: PAGE <= 12'd312;
            12'd997: PAGE <= 12'd834;
            12'd998: PAGE <= 12'd1356;
            12'd999: PAGE <= 12'd1878;
            12'd1000: PAGE <= 12'd347;
            12'd1001: PAGE <= 12'd869;
            12'd1002: PAGE <= 12'd1391;
            12'd1003: PAGE <= 12'd1913;
            12'd1004: PAGE <= 12'd382;
            12'd1005: PAGE <= 12'd904;
            12'd1006: PAGE <= 12'd1426;
            12'd1007: PAGE <= 12'd1948;
            12'd1008: PAGE <= 12'd417;
            12'd1009: PAGE <= 12'd939;
            12'd1010: PAGE <= 12'd1461;
            12'd1011: PAGE <= 12'd1983;
            12'd1012: PAGE <= 12'd452;
            12'd1013: PAGE <= 12'd974;
            12'd1014: PAGE <= 12'd1496;
            12'd1015: PAGE <= 12'd2018;
            12'd1016: PAGE <= 12'd487;
            12'd1017: PAGE <= 12'd1009;
            12'd1018: PAGE <= 12'd1531;
            12'd1019: PAGE <= 12'd0;
            12'd1020: PAGE <= 12'd522;
            12'd1021: PAGE <= 12'd1044;
            12'd1022: PAGE <= 12'd1566;
            12'd1023: PAGE <= 12'd35;
            12'd1024: PAGE <= 12'd557;
            12'd1025: PAGE <= 12'd1079;
            12'd1026: PAGE <= 12'd1601;
            12'd1027: PAGE <= 12'd70;
            12'd1028: PAGE <= 12'd592;
            12'd1029: PAGE <= 12'd1114;
            12'd1030: PAGE <= 12'd1636;
            12'd1031: PAGE <= 12'd105;
            12'd1032: PAGE <= 12'd627;
            12'd1033: PAGE <= 12'd1149;
            12'd1034: PAGE <= 12'd1671;
            12'd1035: PAGE <= 12'd140;
            12'd1036: PAGE <= 12'd662;
            12'd1037: PAGE <= 12'd1184;
            12'd1038: PAGE <= 12'd1706;
            12'd1039: PAGE <= 12'd175;
            12'd1040: PAGE <= 12'd697;
            12'd1041: PAGE <= 12'd1219;
            12'd1042: PAGE <= 12'd1741;
            12'd1043: PAGE <= 12'd210;
            12'd1044: PAGE <= 12'd732;
            12'd1045: PAGE <= 12'd1254;
            12'd1046: PAGE <= 12'd1776;
            12'd1047: PAGE <= 12'd245;
            12'd1048: PAGE <= 12'd767;
            12'd1049: PAGE <= 12'd1289;
            12'd1050: PAGE <= 12'd1811;
            12'd1051: PAGE <= 12'd280;
            12'd1052: PAGE <= 12'd802;
            12'd1053: PAGE <= 12'd1324;
            12'd1054: PAGE <= 12'd1846;
            12'd1055: PAGE <= 12'd315;
            12'd1056: PAGE <= 12'd837;
            12'd1057: PAGE <= 12'd1359;
            12'd1058: PAGE <= 12'd1881;
            12'd1059: PAGE <= 12'd350;
            12'd1060: PAGE <= 12'd872;
            12'd1061: PAGE <= 12'd1394;
            12'd1062: PAGE <= 12'd1916;
            12'd1063: PAGE <= 12'd385;
            12'd1064: PAGE <= 12'd907;
            12'd1065: PAGE <= 12'd1429;
            12'd1066: PAGE <= 12'd1951;
            12'd1067: PAGE <= 12'd420;
            12'd1068: PAGE <= 12'd942;
            12'd1069: PAGE <= 12'd1464;
            12'd1070: PAGE <= 12'd1986;
            12'd1071: PAGE <= 12'd455;
            12'd1072: PAGE <= 12'd977;
            12'd1073: PAGE <= 12'd1499;
            12'd1074: PAGE <= 12'd2021;
            12'd1075: PAGE <= 12'd490;
            12'd1076: PAGE <= 12'd1012;
            12'd1077: PAGE <= 12'd1534;
            12'd1078: PAGE <= 12'd3;
            12'd1079: PAGE <= 12'd525;
            12'd1080: PAGE <= 12'd1047;
            12'd1081: PAGE <= 12'd1569;
            12'd1082: PAGE <= 12'd38;
            12'd1083: PAGE <= 12'd560;
            12'd1084: PAGE <= 12'd1082;
            12'd1085: PAGE <= 12'd1604;
            12'd1086: PAGE <= 12'd73;
            12'd1087: PAGE <= 12'd595;
            12'd1088: PAGE <= 12'd1117;
            12'd1089: PAGE <= 12'd1639;
            12'd1090: PAGE <= 12'd108;
            12'd1091: PAGE <= 12'd630;
            12'd1092: PAGE <= 12'd1152;
            12'd1093: PAGE <= 12'd1674;
            12'd1094: PAGE <= 12'd143;
            12'd1095: PAGE <= 12'd665;
            12'd1096: PAGE <= 12'd1187;
            12'd1097: PAGE <= 12'd1709;
            12'd1098: PAGE <= 12'd178;
            12'd1099: PAGE <= 12'd700;
            12'd1100: PAGE <= 12'd1222;
            12'd1101: PAGE <= 12'd1744;
            12'd1102: PAGE <= 12'd213;
            12'd1103: PAGE <= 12'd735;
            12'd1104: PAGE <= 12'd1257;
            12'd1105: PAGE <= 12'd1779;
            12'd1106: PAGE <= 12'd248;
            12'd1107: PAGE <= 12'd770;
            12'd1108: PAGE <= 12'd1292;
            12'd1109: PAGE <= 12'd1814;
            12'd1110: PAGE <= 12'd283;
            12'd1111: PAGE <= 12'd805;
            12'd1112: PAGE <= 12'd1327;
            12'd1113: PAGE <= 12'd1849;
            12'd1114: PAGE <= 12'd318;
            12'd1115: PAGE <= 12'd840;
            12'd1116: PAGE <= 12'd1362;
            12'd1117: PAGE <= 12'd1884;
            12'd1118: PAGE <= 12'd353;
            12'd1119: PAGE <= 12'd875;
            12'd1120: PAGE <= 12'd1397;
            12'd1121: PAGE <= 12'd1919;
            12'd1122: PAGE <= 12'd388;
            12'd1123: PAGE <= 12'd910;
            12'd1124: PAGE <= 12'd1432;
            12'd1125: PAGE <= 12'd1954;
            12'd1126: PAGE <= 12'd423;
            12'd1127: PAGE <= 12'd945;
            12'd1128: PAGE <= 12'd1467;
            12'd1129: PAGE <= 12'd1989;
            12'd1130: PAGE <= 12'd458;
            12'd1131: PAGE <= 12'd980;
            12'd1132: PAGE <= 12'd1502;
            12'd1133: PAGE <= 12'd2024;
            12'd1134: PAGE <= 12'd493;
            12'd1135: PAGE <= 12'd1015;
            12'd1136: PAGE <= 12'd1537;
            12'd1137: PAGE <= 12'd6;
            12'd1138: PAGE <= 12'd528;
            12'd1139: PAGE <= 12'd1050;
            12'd1140: PAGE <= 12'd1572;
            12'd1141: PAGE <= 12'd41;
            12'd1142: PAGE <= 12'd563;
            12'd1143: PAGE <= 12'd1085;
            12'd1144: PAGE <= 12'd1607;
            12'd1145: PAGE <= 12'd76;
            12'd1146: PAGE <= 12'd598;
            12'd1147: PAGE <= 12'd1120;
            12'd1148: PAGE <= 12'd1642;
            12'd1149: PAGE <= 12'd111;
            12'd1150: PAGE <= 12'd633;
            12'd1151: PAGE <= 12'd1155;
            12'd1152: PAGE <= 12'd1677;
            12'd1153: PAGE <= 12'd146;
            12'd1154: PAGE <= 12'd668;
            12'd1155: PAGE <= 12'd1190;
            12'd1156: PAGE <= 12'd1712;
            12'd1157: PAGE <= 12'd181;
            12'd1158: PAGE <= 12'd703;
            12'd1159: PAGE <= 12'd1225;
            12'd1160: PAGE <= 12'd1747;
            12'd1161: PAGE <= 12'd216;
            12'd1162: PAGE <= 12'd738;
            12'd1163: PAGE <= 12'd1260;
            12'd1164: PAGE <= 12'd1782;
            12'd1165: PAGE <= 12'd251;
            12'd1166: PAGE <= 12'd773;
            12'd1167: PAGE <= 12'd1295;
            12'd1168: PAGE <= 12'd1817;
            12'd1169: PAGE <= 12'd286;
            12'd1170: PAGE <= 12'd808;
            12'd1171: PAGE <= 12'd1330;
            12'd1172: PAGE <= 12'd1852;
            12'd1173: PAGE <= 12'd321;
            12'd1174: PAGE <= 12'd843;
            12'd1175: PAGE <= 12'd1365;
            12'd1176: PAGE <= 12'd1887;
            12'd1177: PAGE <= 12'd356;
            12'd1178: PAGE <= 12'd878;
            12'd1179: PAGE <= 12'd1400;
            12'd1180: PAGE <= 12'd1922;
            12'd1181: PAGE <= 12'd391;
            12'd1182: PAGE <= 12'd913;
            12'd1183: PAGE <= 12'd1435;
            12'd1184: PAGE <= 12'd1957;
            12'd1185: PAGE <= 12'd426;
            12'd1186: PAGE <= 12'd948;
            12'd1187: PAGE <= 12'd1470;
            12'd1188: PAGE <= 12'd1992;
            12'd1189: PAGE <= 12'd461;
            12'd1190: PAGE <= 12'd983;
            12'd1191: PAGE <= 12'd1505;
            12'd1192: PAGE <= 12'd2027;
            12'd1193: PAGE <= 12'd496;
            12'd1194: PAGE <= 12'd1018;
            12'd1195: PAGE <= 12'd1540;
            12'd1196: PAGE <= 12'd9;
            12'd1197: PAGE <= 12'd531;
            12'd1198: PAGE <= 12'd1053;
            12'd1199: PAGE <= 12'd1575;
            12'd1200: PAGE <= 12'd44;
            12'd1201: PAGE <= 12'd566;
            12'd1202: PAGE <= 12'd1088;
            12'd1203: PAGE <= 12'd1610;
            12'd1204: PAGE <= 12'd79;
            12'd1205: PAGE <= 12'd601;
            12'd1206: PAGE <= 12'd1123;
            12'd1207: PAGE <= 12'd1645;
            12'd1208: PAGE <= 12'd114;
            12'd1209: PAGE <= 12'd636;
            12'd1210: PAGE <= 12'd1158;
            12'd1211: PAGE <= 12'd1680;
            12'd1212: PAGE <= 12'd149;
            12'd1213: PAGE <= 12'd671;
            12'd1214: PAGE <= 12'd1193;
            12'd1215: PAGE <= 12'd1715;
            12'd1216: PAGE <= 12'd184;
            12'd1217: PAGE <= 12'd706;
            12'd1218: PAGE <= 12'd1228;
            12'd1219: PAGE <= 12'd1750;
            12'd1220: PAGE <= 12'd219;
            12'd1221: PAGE <= 12'd741;
            12'd1222: PAGE <= 12'd1263;
            12'd1223: PAGE <= 12'd1785;
            12'd1224: PAGE <= 12'd254;
            12'd1225: PAGE <= 12'd776;
            12'd1226: PAGE <= 12'd1298;
            12'd1227: PAGE <= 12'd1820;
            12'd1228: PAGE <= 12'd289;
            12'd1229: PAGE <= 12'd811;
            12'd1230: PAGE <= 12'd1333;
            12'd1231: PAGE <= 12'd1855;
            12'd1232: PAGE <= 12'd324;
            12'd1233: PAGE <= 12'd846;
            12'd1234: PAGE <= 12'd1368;
            12'd1235: PAGE <= 12'd1890;
            12'd1236: PAGE <= 12'd359;
            12'd1237: PAGE <= 12'd881;
            12'd1238: PAGE <= 12'd1403;
            12'd1239: PAGE <= 12'd1925;
            12'd1240: PAGE <= 12'd394;
            12'd1241: PAGE <= 12'd916;
            12'd1242: PAGE <= 12'd1438;
            12'd1243: PAGE <= 12'd1960;
            12'd1244: PAGE <= 12'd429;
            12'd1245: PAGE <= 12'd951;
            12'd1246: PAGE <= 12'd1473;
            12'd1247: PAGE <= 12'd1995;
            12'd1248: PAGE <= 12'd464;
            12'd1249: PAGE <= 12'd986;
            12'd1250: PAGE <= 12'd1508;
            12'd1251: PAGE <= 12'd2030;
            12'd1252: PAGE <= 12'd499;
            12'd1253: PAGE <= 12'd1021;
            12'd1254: PAGE <= 12'd1543;
            12'd1255: PAGE <= 12'd12;
            12'd1256: PAGE <= 12'd534;
            12'd1257: PAGE <= 12'd1056;
            12'd1258: PAGE <= 12'd1578;
            12'd1259: PAGE <= 12'd47;
            12'd1260: PAGE <= 12'd569;
            12'd1261: PAGE <= 12'd1091;
            12'd1262: PAGE <= 12'd1613;
            12'd1263: PAGE <= 12'd82;
            12'd1264: PAGE <= 12'd604;
            12'd1265: PAGE <= 12'd1126;
            12'd1266: PAGE <= 12'd1648;
            12'd1267: PAGE <= 12'd117;
            12'd1268: PAGE <= 12'd639;
            12'd1269: PAGE <= 12'd1161;
            12'd1270: PAGE <= 12'd1683;
            12'd1271: PAGE <= 12'd152;
            12'd1272: PAGE <= 12'd674;
            12'd1273: PAGE <= 12'd1196;
            12'd1274: PAGE <= 12'd1718;
            12'd1275: PAGE <= 12'd187;
            12'd1276: PAGE <= 12'd709;
            12'd1277: PAGE <= 12'd1231;
            12'd1278: PAGE <= 12'd1753;
            12'd1279: PAGE <= 12'd222;
            12'd1280: PAGE <= 12'd744;
            12'd1281: PAGE <= 12'd1266;
            12'd1282: PAGE <= 12'd1788;
            12'd1283: PAGE <= 12'd257;
            12'd1284: PAGE <= 12'd779;
            12'd1285: PAGE <= 12'd1301;
            12'd1286: PAGE <= 12'd1823;
            12'd1287: PAGE <= 12'd292;
            12'd1288: PAGE <= 12'd814;
            12'd1289: PAGE <= 12'd1336;
            12'd1290: PAGE <= 12'd1858;
            12'd1291: PAGE <= 12'd327;
            12'd1292: PAGE <= 12'd849;
            12'd1293: PAGE <= 12'd1371;
            12'd1294: PAGE <= 12'd1893;
            12'd1295: PAGE <= 12'd362;
            12'd1296: PAGE <= 12'd884;
            12'd1297: PAGE <= 12'd1406;
            12'd1298: PAGE <= 12'd1928;
            12'd1299: PAGE <= 12'd397;
            12'd1300: PAGE <= 12'd919;
            12'd1301: PAGE <= 12'd1441;
            12'd1302: PAGE <= 12'd1963;
            12'd1303: PAGE <= 12'd432;
            12'd1304: PAGE <= 12'd954;
            12'd1305: PAGE <= 12'd1476;
            12'd1306: PAGE <= 12'd1998;
            12'd1307: PAGE <= 12'd467;
            12'd1308: PAGE <= 12'd989;
            12'd1309: PAGE <= 12'd1511;
            12'd1310: PAGE <= 12'd2033;
            12'd1311: PAGE <= 12'd502;
            12'd1312: PAGE <= 12'd1024;
            12'd1313: PAGE <= 12'd1546;
            12'd1314: PAGE <= 12'd15;
            12'd1315: PAGE <= 12'd537;
            12'd1316: PAGE <= 12'd1059;
            12'd1317: PAGE <= 12'd1581;
            12'd1318: PAGE <= 12'd50;
            12'd1319: PAGE <= 12'd572;
            12'd1320: PAGE <= 12'd1094;
            12'd1321: PAGE <= 12'd1616;
            12'd1322: PAGE <= 12'd85;
            12'd1323: PAGE <= 12'd607;
            12'd1324: PAGE <= 12'd1129;
            12'd1325: PAGE <= 12'd1651;
            12'd1326: PAGE <= 12'd120;
            12'd1327: PAGE <= 12'd642;
            12'd1328: PAGE <= 12'd1164;
            12'd1329: PAGE <= 12'd1686;
            12'd1330: PAGE <= 12'd155;
            12'd1331: PAGE <= 12'd677;
            12'd1332: PAGE <= 12'd1199;
            12'd1333: PAGE <= 12'd1721;
            12'd1334: PAGE <= 12'd190;
            12'd1335: PAGE <= 12'd712;
            12'd1336: PAGE <= 12'd1234;
            12'd1337: PAGE <= 12'd1756;
            12'd1338: PAGE <= 12'd225;
            12'd1339: PAGE <= 12'd747;
            12'd1340: PAGE <= 12'd1269;
            12'd1341: PAGE <= 12'd1791;
            12'd1342: PAGE <= 12'd260;
            12'd1343: PAGE <= 12'd782;
            12'd1344: PAGE <= 12'd1304;
            12'd1345: PAGE <= 12'd1826;
            12'd1346: PAGE <= 12'd295;
            12'd1347: PAGE <= 12'd817;
            12'd1348: PAGE <= 12'd1339;
            12'd1349: PAGE <= 12'd1861;
            12'd1350: PAGE <= 12'd330;
            12'd1351: PAGE <= 12'd852;
            12'd1352: PAGE <= 12'd1374;
            12'd1353: PAGE <= 12'd1896;
            12'd1354: PAGE <= 12'd365;
            12'd1355: PAGE <= 12'd887;
            12'd1356: PAGE <= 12'd1409;
            12'd1357: PAGE <= 12'd1931;
            12'd1358: PAGE <= 12'd400;
            12'd1359: PAGE <= 12'd922;
            12'd1360: PAGE <= 12'd1444;
            12'd1361: PAGE <= 12'd1966;
            12'd1362: PAGE <= 12'd435;
            12'd1363: PAGE <= 12'd957;
            12'd1364: PAGE <= 12'd1479;
            12'd1365: PAGE <= 12'd2001;
            12'd1366: PAGE <= 12'd470;
            12'd1367: PAGE <= 12'd992;
            12'd1368: PAGE <= 12'd1514;
            12'd1369: PAGE <= 12'd2036;
            12'd1370: PAGE <= 12'd505;
            12'd1371: PAGE <= 12'd1027;
            12'd1372: PAGE <= 12'd1549;
            12'd1373: PAGE <= 12'd18;
            12'd1374: PAGE <= 12'd540;
            12'd1375: PAGE <= 12'd1062;
            12'd1376: PAGE <= 12'd1584;
            12'd1377: PAGE <= 12'd53;
            12'd1378: PAGE <= 12'd575;
            12'd1379: PAGE <= 12'd1097;
            12'd1380: PAGE <= 12'd1619;
            12'd1381: PAGE <= 12'd88;
            12'd1382: PAGE <= 12'd610;
            12'd1383: PAGE <= 12'd1132;
            12'd1384: PAGE <= 12'd1654;
            12'd1385: PAGE <= 12'd123;
            12'd1386: PAGE <= 12'd645;
            12'd1387: PAGE <= 12'd1167;
            12'd1388: PAGE <= 12'd1689;
            12'd1389: PAGE <= 12'd158;
            12'd1390: PAGE <= 12'd680;
            12'd1391: PAGE <= 12'd1202;
            12'd1392: PAGE <= 12'd1724;
            12'd1393: PAGE <= 12'd193;
            12'd1394: PAGE <= 12'd715;
            12'd1395: PAGE <= 12'd1237;
            12'd1396: PAGE <= 12'd1759;
            12'd1397: PAGE <= 12'd228;
            12'd1398: PAGE <= 12'd750;
            12'd1399: PAGE <= 12'd1272;
            12'd1400: PAGE <= 12'd1794;
            12'd1401: PAGE <= 12'd263;
            12'd1402: PAGE <= 12'd785;
            12'd1403: PAGE <= 12'd1307;
            12'd1404: PAGE <= 12'd1829;
            12'd1405: PAGE <= 12'd298;
            12'd1406: PAGE <= 12'd820;
            12'd1407: PAGE <= 12'd1342;
            12'd1408: PAGE <= 12'd1864;
            12'd1409: PAGE <= 12'd333;
            12'd1410: PAGE <= 12'd855;
            12'd1411: PAGE <= 12'd1377;
            12'd1412: PAGE <= 12'd1899;
            12'd1413: PAGE <= 12'd368;
            12'd1414: PAGE <= 12'd890;
            12'd1415: PAGE <= 12'd1412;
            12'd1416: PAGE <= 12'd1934;
            12'd1417: PAGE <= 12'd403;
            12'd1418: PAGE <= 12'd925;
            12'd1419: PAGE <= 12'd1447;
            12'd1420: PAGE <= 12'd1969;
            12'd1421: PAGE <= 12'd438;
            12'd1422: PAGE <= 12'd960;
            12'd1423: PAGE <= 12'd1482;
            12'd1424: PAGE <= 12'd2004;
            12'd1425: PAGE <= 12'd473;
            12'd1426: PAGE <= 12'd995;
            12'd1427: PAGE <= 12'd1517;
            12'd1428: PAGE <= 12'd2039;
            12'd1429: PAGE <= 12'd508;
            12'd1430: PAGE <= 12'd1030;
            12'd1431: PAGE <= 12'd1552;
            12'd1432: PAGE <= 12'd21;
            12'd1433: PAGE <= 12'd543;
            12'd1434: PAGE <= 12'd1065;
            12'd1435: PAGE <= 12'd1587;
            12'd1436: PAGE <= 12'd56;
            12'd1437: PAGE <= 12'd578;
            12'd1438: PAGE <= 12'd1100;
            12'd1439: PAGE <= 12'd1622;
            12'd1440: PAGE <= 12'd91;
            12'd1441: PAGE <= 12'd613;
            12'd1442: PAGE <= 12'd1135;
            12'd1443: PAGE <= 12'd1657;
            12'd1444: PAGE <= 12'd126;
            12'd1445: PAGE <= 12'd648;
            12'd1446: PAGE <= 12'd1170;
            12'd1447: PAGE <= 12'd1692;
            12'd1448: PAGE <= 12'd161;
            12'd1449: PAGE <= 12'd683;
            12'd1450: PAGE <= 12'd1205;
            12'd1451: PAGE <= 12'd1727;
            12'd1452: PAGE <= 12'd196;
            12'd1453: PAGE <= 12'd718;
            12'd1454: PAGE <= 12'd1240;
            12'd1455: PAGE <= 12'd1762;
            12'd1456: PAGE <= 12'd231;
            12'd1457: PAGE <= 12'd753;
            12'd1458: PAGE <= 12'd1275;
            12'd1459: PAGE <= 12'd1797;
            12'd1460: PAGE <= 12'd266;
            12'd1461: PAGE <= 12'd788;
            12'd1462: PAGE <= 12'd1310;
            12'd1463: PAGE <= 12'd1832;
            12'd1464: PAGE <= 12'd301;
            12'd1465: PAGE <= 12'd823;
            12'd1466: PAGE <= 12'd1345;
            12'd1467: PAGE <= 12'd1867;
            12'd1468: PAGE <= 12'd336;
            12'd1469: PAGE <= 12'd858;
            12'd1470: PAGE <= 12'd1380;
            12'd1471: PAGE <= 12'd1902;
            12'd1472: PAGE <= 12'd371;
            12'd1473: PAGE <= 12'd893;
            12'd1474: PAGE <= 12'd1415;
            12'd1475: PAGE <= 12'd1937;
            12'd1476: PAGE <= 12'd406;
            12'd1477: PAGE <= 12'd928;
            12'd1478: PAGE <= 12'd1450;
            12'd1479: PAGE <= 12'd1972;
            12'd1480: PAGE <= 12'd441;
            12'd1481: PAGE <= 12'd963;
            12'd1482: PAGE <= 12'd1485;
            12'd1483: PAGE <= 12'd2007;
            12'd1484: PAGE <= 12'd476;
            12'd1485: PAGE <= 12'd998;
            12'd1486: PAGE <= 12'd1520;
            12'd1487: PAGE <= 12'd2042;
            12'd1488: PAGE <= 12'd511;
            12'd1489: PAGE <= 12'd1033;
            12'd1490: PAGE <= 12'd1555;
            12'd1491: PAGE <= 12'd24;
            12'd1492: PAGE <= 12'd546;
            12'd1493: PAGE <= 12'd1068;
            12'd1494: PAGE <= 12'd1590;
            12'd1495: PAGE <= 12'd59;
            12'd1496: PAGE <= 12'd581;
            12'd1497: PAGE <= 12'd1103;
            12'd1498: PAGE <= 12'd1625;
            12'd1499: PAGE <= 12'd94;
            12'd1500: PAGE <= 12'd616;
            12'd1501: PAGE <= 12'd1138;
            12'd1502: PAGE <= 12'd1660;
            12'd1503: PAGE <= 12'd129;
            12'd1504: PAGE <= 12'd651;
            12'd1505: PAGE <= 12'd1173;
            12'd1506: PAGE <= 12'd1695;
            12'd1507: PAGE <= 12'd164;
            12'd1508: PAGE <= 12'd686;
            12'd1509: PAGE <= 12'd1208;
            12'd1510: PAGE <= 12'd1730;
            12'd1511: PAGE <= 12'd199;
            12'd1512: PAGE <= 12'd721;
            12'd1513: PAGE <= 12'd1243;
            12'd1514: PAGE <= 12'd1765;
            12'd1515: PAGE <= 12'd234;
            12'd1516: PAGE <= 12'd756;
            12'd1517: PAGE <= 12'd1278;
            12'd1518: PAGE <= 12'd1800;
            12'd1519: PAGE <= 12'd269;
            12'd1520: PAGE <= 12'd791;
            12'd1521: PAGE <= 12'd1313;
            12'd1522: PAGE <= 12'd1835;
            12'd1523: PAGE <= 12'd304;
            12'd1524: PAGE <= 12'd826;
            12'd1525: PAGE <= 12'd1348;
            12'd1526: PAGE <= 12'd1870;
            12'd1527: PAGE <= 12'd339;
            12'd1528: PAGE <= 12'd861;
            12'd1529: PAGE <= 12'd1383;
            12'd1530: PAGE <= 12'd1905;
            12'd1531: PAGE <= 12'd374;
            12'd1532: PAGE <= 12'd896;
            12'd1533: PAGE <= 12'd1418;
            12'd1534: PAGE <= 12'd1940;
            12'd1535: PAGE <= 12'd409;
            12'd1536: PAGE <= 12'd931;
            12'd1537: PAGE <= 12'd1453;
            12'd1538: PAGE <= 12'd1975;
            12'd1539: PAGE <= 12'd444;
            12'd1540: PAGE <= 12'd966;
            12'd1541: PAGE <= 12'd1488;
            12'd1542: PAGE <= 12'd2010;
            12'd1543: PAGE <= 12'd479;
            12'd1544: PAGE <= 12'd1001;
            12'd1545: PAGE <= 12'd1523;
            12'd1546: PAGE <= 12'd2045;
            12'd1547: PAGE <= 12'd514;
            12'd1548: PAGE <= 12'd1036;
            12'd1549: PAGE <= 12'd1558;
            12'd1550: PAGE <= 12'd27;
            12'd1551: PAGE <= 12'd549;
            12'd1552: PAGE <= 12'd1071;
            12'd1553: PAGE <= 12'd1593;
            12'd1554: PAGE <= 12'd62;
            12'd1555: PAGE <= 12'd584;
            12'd1556: PAGE <= 12'd1106;
            12'd1557: PAGE <= 12'd1628;
            12'd1558: PAGE <= 12'd97;
            12'd1559: PAGE <= 12'd619;
            12'd1560: PAGE <= 12'd1141;
            12'd1561: PAGE <= 12'd1663;
            12'd1562: PAGE <= 12'd132;
            12'd1563: PAGE <= 12'd654;
            12'd1564: PAGE <= 12'd1176;
            12'd1565: PAGE <= 12'd1698;
            12'd1566: PAGE <= 12'd167;
            12'd1567: PAGE <= 12'd689;
            12'd1568: PAGE <= 12'd1211;
            12'd1569: PAGE <= 12'd1733;
            12'd1570: PAGE <= 12'd202;
            12'd1571: PAGE <= 12'd724;
            12'd1572: PAGE <= 12'd1246;
            12'd1573: PAGE <= 12'd1768;
            12'd1574: PAGE <= 12'd237;
            12'd1575: PAGE <= 12'd759;
            12'd1576: PAGE <= 12'd1281;
            12'd1577: PAGE <= 12'd1803;
            12'd1578: PAGE <= 12'd272;
            12'd1579: PAGE <= 12'd794;
            12'd1580: PAGE <= 12'd1316;
            12'd1581: PAGE <= 12'd1838;
            12'd1582: PAGE <= 12'd307;
            12'd1583: PAGE <= 12'd829;
            12'd1584: PAGE <= 12'd1351;
            12'd1585: PAGE <= 12'd1873;
            12'd1586: PAGE <= 12'd342;
            12'd1587: PAGE <= 12'd864;
            12'd1588: PAGE <= 12'd1386;
            12'd1589: PAGE <= 12'd1908;
            12'd1590: PAGE <= 12'd377;
            12'd1591: PAGE <= 12'd899;
            12'd1592: PAGE <= 12'd1421;
            12'd1593: PAGE <= 12'd1943;
            12'd1594: PAGE <= 12'd412;
            12'd1595: PAGE <= 12'd934;
            12'd1596: PAGE <= 12'd1456;
            12'd1597: PAGE <= 12'd1978;
            12'd1598: PAGE <= 12'd447;
            12'd1599: PAGE <= 12'd969;
            12'd1600: PAGE <= 12'd1491;
            12'd1601: PAGE <= 12'd2013;
            12'd1602: PAGE <= 12'd482;
            12'd1603: PAGE <= 12'd1004;
            12'd1604: PAGE <= 12'd1526;
            12'd1605: PAGE <= 12'd2048;
            12'd1606: PAGE <= 12'd517;
            12'd1607: PAGE <= 12'd1039;
            12'd1608: PAGE <= 12'd1561;
            12'd1609: PAGE <= 12'd30;
            12'd1610: PAGE <= 12'd552;
            12'd1611: PAGE <= 12'd1074;
            12'd1612: PAGE <= 12'd1596;
            12'd1613: PAGE <= 12'd65;
            12'd1614: PAGE <= 12'd587;
            12'd1615: PAGE <= 12'd1109;
            12'd1616: PAGE <= 12'd1631;
            12'd1617: PAGE <= 12'd100;
            12'd1618: PAGE <= 12'd622;
            12'd1619: PAGE <= 12'd1144;
            12'd1620: PAGE <= 12'd1666;
            12'd1621: PAGE <= 12'd135;
            12'd1622: PAGE <= 12'd657;
            12'd1623: PAGE <= 12'd1179;
            12'd1624: PAGE <= 12'd1701;
            12'd1625: PAGE <= 12'd170;
            12'd1626: PAGE <= 12'd692;
            12'd1627: PAGE <= 12'd1214;
            12'd1628: PAGE <= 12'd1736;
            12'd1629: PAGE <= 12'd205;
            12'd1630: PAGE <= 12'd727;
            12'd1631: PAGE <= 12'd1249;
            12'd1632: PAGE <= 12'd1771;
            12'd1633: PAGE <= 12'd240;
            12'd1634: PAGE <= 12'd762;
            12'd1635: PAGE <= 12'd1284;
            12'd1636: PAGE <= 12'd1806;
            12'd1637: PAGE <= 12'd275;
            12'd1638: PAGE <= 12'd797;
            12'd1639: PAGE <= 12'd1319;
            12'd1640: PAGE <= 12'd1841;
            12'd1641: PAGE <= 12'd310;
            12'd1642: PAGE <= 12'd832;
            12'd1643: PAGE <= 12'd1354;
            12'd1644: PAGE <= 12'd1876;
            12'd1645: PAGE <= 12'd345;
            12'd1646: PAGE <= 12'd867;
            12'd1647: PAGE <= 12'd1389;
            12'd1648: PAGE <= 12'd1911;
            12'd1649: PAGE <= 12'd380;
            12'd1650: PAGE <= 12'd902;
            12'd1651: PAGE <= 12'd1424;
            12'd1652: PAGE <= 12'd1946;
            12'd1653: PAGE <= 12'd415;
            12'd1654: PAGE <= 12'd937;
            12'd1655: PAGE <= 12'd1459;
            12'd1656: PAGE <= 12'd1981;
            12'd1657: PAGE <= 12'd450;
            12'd1658: PAGE <= 12'd972;
            12'd1659: PAGE <= 12'd1494;
            12'd1660: PAGE <= 12'd2016;
            12'd1661: PAGE <= 12'd485;
            12'd1662: PAGE <= 12'd1007;
            12'd1663: PAGE <= 12'd1529;
            12'd1664: PAGE <= 12'd2051;
            12'd1665: PAGE <= 12'd520;
            12'd1666: PAGE <= 12'd1042;
            12'd1667: PAGE <= 12'd1564;
            12'd1668: PAGE <= 12'd33;
            12'd1669: PAGE <= 12'd555;
            12'd1670: PAGE <= 12'd1077;
            12'd1671: PAGE <= 12'd1599;
            12'd1672: PAGE <= 12'd68;
            12'd1673: PAGE <= 12'd590;
            12'd1674: PAGE <= 12'd1112;
            12'd1675: PAGE <= 12'd1634;
            12'd1676: PAGE <= 12'd103;
            12'd1677: PAGE <= 12'd625;
            12'd1678: PAGE <= 12'd1147;
            12'd1679: PAGE <= 12'd1669;
            12'd1680: PAGE <= 12'd138;
            12'd1681: PAGE <= 12'd660;
            12'd1682: PAGE <= 12'd1182;
            12'd1683: PAGE <= 12'd1704;
            12'd1684: PAGE <= 12'd173;
            12'd1685: PAGE <= 12'd695;
            12'd1686: PAGE <= 12'd1217;
            12'd1687: PAGE <= 12'd1739;
            12'd1688: PAGE <= 12'd208;
            12'd1689: PAGE <= 12'd730;
            12'd1690: PAGE <= 12'd1252;
            12'd1691: PAGE <= 12'd1774;
            12'd1692: PAGE <= 12'd243;
            12'd1693: PAGE <= 12'd765;
            12'd1694: PAGE <= 12'd1287;
            12'd1695: PAGE <= 12'd1809;
            12'd1696: PAGE <= 12'd278;
            12'd1697: PAGE <= 12'd800;
            12'd1698: PAGE <= 12'd1322;
            12'd1699: PAGE <= 12'd1844;
            12'd1700: PAGE <= 12'd313;
            12'd1701: PAGE <= 12'd835;
            12'd1702: PAGE <= 12'd1357;
            12'd1703: PAGE <= 12'd1879;
            12'd1704: PAGE <= 12'd348;
            12'd1705: PAGE <= 12'd870;
            12'd1706: PAGE <= 12'd1392;
            12'd1707: PAGE <= 12'd1914;
            12'd1708: PAGE <= 12'd383;
            12'd1709: PAGE <= 12'd905;
            12'd1710: PAGE <= 12'd1427;
            12'd1711: PAGE <= 12'd1949;
            12'd1712: PAGE <= 12'd418;
            12'd1713: PAGE <= 12'd940;
            12'd1714: PAGE <= 12'd1462;
            12'd1715: PAGE <= 12'd1984;
            12'd1716: PAGE <= 12'd453;
            12'd1717: PAGE <= 12'd975;
            12'd1718: PAGE <= 12'd1497;
            12'd1719: PAGE <= 12'd2019;
            12'd1720: PAGE <= 12'd488;
            12'd1721: PAGE <= 12'd1010;
            12'd1722: PAGE <= 12'd1532;
            12'd1723: PAGE <= 12'd1;
            12'd1724: PAGE <= 12'd523;
            12'd1725: PAGE <= 12'd1045;
            12'd1726: PAGE <= 12'd1567;
            12'd1727: PAGE <= 12'd36;
            12'd1728: PAGE <= 12'd558;
            12'd1729: PAGE <= 12'd1080;
            12'd1730: PAGE <= 12'd1602;
            12'd1731: PAGE <= 12'd71;
            12'd1732: PAGE <= 12'd593;
            12'd1733: PAGE <= 12'd1115;
            12'd1734: PAGE <= 12'd1637;
            12'd1735: PAGE <= 12'd106;
            12'd1736: PAGE <= 12'd628;
            12'd1737: PAGE <= 12'd1150;
            12'd1738: PAGE <= 12'd1672;
            12'd1739: PAGE <= 12'd141;
            12'd1740: PAGE <= 12'd663;
            12'd1741: PAGE <= 12'd1185;
            12'd1742: PAGE <= 12'd1707;
            12'd1743: PAGE <= 12'd176;
            12'd1744: PAGE <= 12'd698;
            12'd1745: PAGE <= 12'd1220;
            12'd1746: PAGE <= 12'd1742;
            12'd1747: PAGE <= 12'd211;
            12'd1748: PAGE <= 12'd733;
            12'd1749: PAGE <= 12'd1255;
            12'd1750: PAGE <= 12'd1777;
            12'd1751: PAGE <= 12'd246;
            12'd1752: PAGE <= 12'd768;
            12'd1753: PAGE <= 12'd1290;
            12'd1754: PAGE <= 12'd1812;
            12'd1755: PAGE <= 12'd281;
            12'd1756: PAGE <= 12'd803;
            12'd1757: PAGE <= 12'd1325;
            12'd1758: PAGE <= 12'd1847;
            12'd1759: PAGE <= 12'd316;
            12'd1760: PAGE <= 12'd838;
            12'd1761: PAGE <= 12'd1360;
            12'd1762: PAGE <= 12'd1882;
            12'd1763: PAGE <= 12'd351;
            12'd1764: PAGE <= 12'd873;
            12'd1765: PAGE <= 12'd1395;
            12'd1766: PAGE <= 12'd1917;
            12'd1767: PAGE <= 12'd386;
            12'd1768: PAGE <= 12'd908;
            12'd1769: PAGE <= 12'd1430;
            12'd1770: PAGE <= 12'd1952;
            12'd1771: PAGE <= 12'd421;
            12'd1772: PAGE <= 12'd943;
            12'd1773: PAGE <= 12'd1465;
            12'd1774: PAGE <= 12'd1987;
            12'd1775: PAGE <= 12'd456;
            12'd1776: PAGE <= 12'd978;
            12'd1777: PAGE <= 12'd1500;
            12'd1778: PAGE <= 12'd2022;
            12'd1779: PAGE <= 12'd491;
            12'd1780: PAGE <= 12'd1013;
            12'd1781: PAGE <= 12'd1535;
            12'd1782: PAGE <= 12'd4;
            12'd1783: PAGE <= 12'd526;
            12'd1784: PAGE <= 12'd1048;
            12'd1785: PAGE <= 12'd1570;
            12'd1786: PAGE <= 12'd39;
            12'd1787: PAGE <= 12'd561;
            12'd1788: PAGE <= 12'd1083;
            12'd1789: PAGE <= 12'd1605;
            12'd1790: PAGE <= 12'd74;
            12'd1791: PAGE <= 12'd596;
            12'd1792: PAGE <= 12'd1118;
            12'd1793: PAGE <= 12'd1640;
            12'd1794: PAGE <= 12'd109;
            12'd1795: PAGE <= 12'd631;
            12'd1796: PAGE <= 12'd1153;
            12'd1797: PAGE <= 12'd1675;
            12'd1798: PAGE <= 12'd144;
            12'd1799: PAGE <= 12'd666;
            12'd1800: PAGE <= 12'd1188;
            12'd1801: PAGE <= 12'd1710;
            12'd1802: PAGE <= 12'd179;
            12'd1803: PAGE <= 12'd701;
            12'd1804: PAGE <= 12'd1223;
            12'd1805: PAGE <= 12'd1745;
            12'd1806: PAGE <= 12'd214;
            12'd1807: PAGE <= 12'd736;
            12'd1808: PAGE <= 12'd1258;
            12'd1809: PAGE <= 12'd1780;
            12'd1810: PAGE <= 12'd249;
            12'd1811: PAGE <= 12'd771;
            12'd1812: PAGE <= 12'd1293;
            12'd1813: PAGE <= 12'd1815;
            12'd1814: PAGE <= 12'd284;
            12'd1815: PAGE <= 12'd806;
            12'd1816: PAGE <= 12'd1328;
            12'd1817: PAGE <= 12'd1850;
            12'd1818: PAGE <= 12'd319;
            12'd1819: PAGE <= 12'd841;
            12'd1820: PAGE <= 12'd1363;
            12'd1821: PAGE <= 12'd1885;
            12'd1822: PAGE <= 12'd354;
            12'd1823: PAGE <= 12'd876;
            12'd1824: PAGE <= 12'd1398;
            12'd1825: PAGE <= 12'd1920;
            12'd1826: PAGE <= 12'd389;
            12'd1827: PAGE <= 12'd911;
            12'd1828: PAGE <= 12'd1433;
            12'd1829: PAGE <= 12'd1955;
            12'd1830: PAGE <= 12'd424;
            12'd1831: PAGE <= 12'd946;
            12'd1832: PAGE <= 12'd1468;
            12'd1833: PAGE <= 12'd1990;
            12'd1834: PAGE <= 12'd459;
            12'd1835: PAGE <= 12'd981;
            12'd1836: PAGE <= 12'd1503;
            12'd1837: PAGE <= 12'd2025;
            12'd1838: PAGE <= 12'd494;
            12'd1839: PAGE <= 12'd1016;
            12'd1840: PAGE <= 12'd1538;
            12'd1841: PAGE <= 12'd7;
            12'd1842: PAGE <= 12'd529;
            12'd1843: PAGE <= 12'd1051;
            12'd1844: PAGE <= 12'd1573;
            12'd1845: PAGE <= 12'd42;
            12'd1846: PAGE <= 12'd564;
            12'd1847: PAGE <= 12'd1086;
            12'd1848: PAGE <= 12'd1608;
            12'd1849: PAGE <= 12'd77;
            12'd1850: PAGE <= 12'd599;
            12'd1851: PAGE <= 12'd1121;
            12'd1852: PAGE <= 12'd1643;
            12'd1853: PAGE <= 12'd112;
            12'd1854: PAGE <= 12'd634;
            12'd1855: PAGE <= 12'd1156;
            12'd1856: PAGE <= 12'd1678;
            12'd1857: PAGE <= 12'd147;
            12'd1858: PAGE <= 12'd669;
            12'd1859: PAGE <= 12'd1191;
            12'd1860: PAGE <= 12'd1713;
            12'd1861: PAGE <= 12'd182;
            12'd1862: PAGE <= 12'd704;
            12'd1863: PAGE <= 12'd1226;
            12'd1864: PAGE <= 12'd1748;
            12'd1865: PAGE <= 12'd217;
            12'd1866: PAGE <= 12'd739;
            12'd1867: PAGE <= 12'd1261;
            12'd1868: PAGE <= 12'd1783;
            12'd1869: PAGE <= 12'd252;
            12'd1870: PAGE <= 12'd774;
            12'd1871: PAGE <= 12'd1296;
            12'd1872: PAGE <= 12'd1818;
            12'd1873: PAGE <= 12'd287;
            12'd1874: PAGE <= 12'd809;
            12'd1875: PAGE <= 12'd1331;
            12'd1876: PAGE <= 12'd1853;
            12'd1877: PAGE <= 12'd322;
            12'd1878: PAGE <= 12'd844;
            12'd1879: PAGE <= 12'd1366;
            12'd1880: PAGE <= 12'd1888;
            12'd1881: PAGE <= 12'd357;
            12'd1882: PAGE <= 12'd879;
            12'd1883: PAGE <= 12'd1401;
            12'd1884: PAGE <= 12'd1923;
            12'd1885: PAGE <= 12'd392;
            12'd1886: PAGE <= 12'd914;
            12'd1887: PAGE <= 12'd1436;
            12'd1888: PAGE <= 12'd1958;
            12'd1889: PAGE <= 12'd427;
            12'd1890: PAGE <= 12'd949;
            12'd1891: PAGE <= 12'd1471;
            12'd1892: PAGE <= 12'd1993;
            12'd1893: PAGE <= 12'd462;
            12'd1894: PAGE <= 12'd984;
            12'd1895: PAGE <= 12'd1506;
            12'd1896: PAGE <= 12'd2028;
            12'd1897: PAGE <= 12'd497;
            12'd1898: PAGE <= 12'd1019;
            12'd1899: PAGE <= 12'd1541;
            12'd1900: PAGE <= 12'd10;
            12'd1901: PAGE <= 12'd532;
            12'd1902: PAGE <= 12'd1054;
            12'd1903: PAGE <= 12'd1576;
            12'd1904: PAGE <= 12'd45;
            12'd1905: PAGE <= 12'd567;
            12'd1906: PAGE <= 12'd1089;
            12'd1907: PAGE <= 12'd1611;
            12'd1908: PAGE <= 12'd80;
            12'd1909: PAGE <= 12'd602;
            12'd1910: PAGE <= 12'd1124;
            12'd1911: PAGE <= 12'd1646;
            12'd1912: PAGE <= 12'd115;
            12'd1913: PAGE <= 12'd637;
            12'd1914: PAGE <= 12'd1159;
            12'd1915: PAGE <= 12'd1681;
            12'd1916: PAGE <= 12'd150;
            12'd1917: PAGE <= 12'd672;
            12'd1918: PAGE <= 12'd1194;
            12'd1919: PAGE <= 12'd1716;
            12'd1920: PAGE <= 12'd185;
            12'd1921: PAGE <= 12'd707;
            12'd1922: PAGE <= 12'd1229;
            12'd1923: PAGE <= 12'd1751;
            12'd1924: PAGE <= 12'd220;
            12'd1925: PAGE <= 12'd742;
            12'd1926: PAGE <= 12'd1264;
            12'd1927: PAGE <= 12'd1786;
            12'd1928: PAGE <= 12'd255;
            12'd1929: PAGE <= 12'd777;
            12'd1930: PAGE <= 12'd1299;
            12'd1931: PAGE <= 12'd1821;
            12'd1932: PAGE <= 12'd290;
            12'd1933: PAGE <= 12'd812;
            12'd1934: PAGE <= 12'd1334;
            12'd1935: PAGE <= 12'd1856;
            12'd1936: PAGE <= 12'd325;
            12'd1937: PAGE <= 12'd847;
            12'd1938: PAGE <= 12'd1369;
            12'd1939: PAGE <= 12'd1891;
            12'd1940: PAGE <= 12'd360;
            12'd1941: PAGE <= 12'd882;
            12'd1942: PAGE <= 12'd1404;
            12'd1943: PAGE <= 12'd1926;
            12'd1944: PAGE <= 12'd395;
            12'd1945: PAGE <= 12'd917;
            12'd1946: PAGE <= 12'd1439;
            12'd1947: PAGE <= 12'd1961;
            12'd1948: PAGE <= 12'd430;
            12'd1949: PAGE <= 12'd952;
            12'd1950: PAGE <= 12'd1474;
            12'd1951: PAGE <= 12'd1996;
            12'd1952: PAGE <= 12'd465;
            12'd1953: PAGE <= 12'd987;
            12'd1954: PAGE <= 12'd1509;
            12'd1955: PAGE <= 12'd2031;
            12'd1956: PAGE <= 12'd500;
            12'd1957: PAGE <= 12'd1022;
            12'd1958: PAGE <= 12'd1544;
            12'd1959: PAGE <= 12'd13;
            12'd1960: PAGE <= 12'd535;
            12'd1961: PAGE <= 12'd1057;
            12'd1962: PAGE <= 12'd1579;
            12'd1963: PAGE <= 12'd48;
            12'd1964: PAGE <= 12'd570;
            12'd1965: PAGE <= 12'd1092;
            12'd1966: PAGE <= 12'd1614;
            12'd1967: PAGE <= 12'd83;
            12'd1968: PAGE <= 12'd605;
            12'd1969: PAGE <= 12'd1127;
            12'd1970: PAGE <= 12'd1649;
            12'd1971: PAGE <= 12'd118;
            12'd1972: PAGE <= 12'd640;
            12'd1973: PAGE <= 12'd1162;
            12'd1974: PAGE <= 12'd1684;
            12'd1975: PAGE <= 12'd153;
            12'd1976: PAGE <= 12'd675;
            12'd1977: PAGE <= 12'd1197;
            12'd1978: PAGE <= 12'd1719;
            12'd1979: PAGE <= 12'd188;
            12'd1980: PAGE <= 12'd710;
            12'd1981: PAGE <= 12'd1232;
            12'd1982: PAGE <= 12'd1754;
            12'd1983: PAGE <= 12'd223;
            12'd1984: PAGE <= 12'd745;
            12'd1985: PAGE <= 12'd1267;
            12'd1986: PAGE <= 12'd1789;
            12'd1987: PAGE <= 12'd258;
            12'd1988: PAGE <= 12'd780;
            12'd1989: PAGE <= 12'd1302;
            12'd1990: PAGE <= 12'd1824;
            12'd1991: PAGE <= 12'd293;
            12'd1992: PAGE <= 12'd815;
            12'd1993: PAGE <= 12'd1337;
            12'd1994: PAGE <= 12'd1859;
            12'd1995: PAGE <= 12'd328;
            12'd1996: PAGE <= 12'd850;
            12'd1997: PAGE <= 12'd1372;
            12'd1998: PAGE <= 12'd1894;
            12'd1999: PAGE <= 12'd363;
            12'd2000: PAGE <= 12'd885;
            12'd2001: PAGE <= 12'd1407;
            12'd2002: PAGE <= 12'd1929;
            12'd2003: PAGE <= 12'd398;
            12'd2004: PAGE <= 12'd920;
            12'd2005: PAGE <= 12'd1442;
            12'd2006: PAGE <= 12'd1964;
            12'd2007: PAGE <= 12'd433;
            12'd2008: PAGE <= 12'd955;
            12'd2009: PAGE <= 12'd1477;
            12'd2010: PAGE <= 12'd1999;
            12'd2011: PAGE <= 12'd468;
            12'd2012: PAGE <= 12'd990;
            12'd2013: PAGE <= 12'd1512;
            12'd2014: PAGE <= 12'd2034;
            12'd2015: PAGE <= 12'd503;
            12'd2016: PAGE <= 12'd1025;
            12'd2017: PAGE <= 12'd1547;
            12'd2018: PAGE <= 12'd16;
            12'd2019: PAGE <= 12'd538;
            12'd2020: PAGE <= 12'd1060;
            12'd2021: PAGE <= 12'd1582;
            12'd2022: PAGE <= 12'd51;
            12'd2023: PAGE <= 12'd573;
            12'd2024: PAGE <= 12'd1095;
            12'd2025: PAGE <= 12'd1617;
            12'd2026: PAGE <= 12'd86;
            12'd2027: PAGE <= 12'd608;
            12'd2028: PAGE <= 12'd1130;
            12'd2029: PAGE <= 12'd1652;
            12'd2030: PAGE <= 12'd121;
            12'd2031: PAGE <= 12'd643;
            12'd2032: PAGE <= 12'd1165;
            12'd2033: PAGE <= 12'd1687;
            12'd2034: PAGE <= 12'd156;
            12'd2035: PAGE <= 12'd678;
            12'd2036: PAGE <= 12'd1200;
            12'd2037: PAGE <= 12'd1722;
            12'd2038: PAGE <= 12'd191;
            12'd2039: PAGE <= 12'd713;
            12'd2040: PAGE <= 12'd1235;
            12'd2041: PAGE <= 12'd1757;
            12'd2042: PAGE <= 12'd226;
            12'd2043: PAGE <= 12'd748;
            12'd2044: PAGE <= 12'd1270;
            12'd2045: PAGE <= 12'd1792;
            12'd2046: PAGE <= 12'd261;
            12'd2047: PAGE <= 12'd783;
            12'd2048: PAGE <= 12'd1305;
            12'd2049: PAGE <= 12'd1827;
            12'd2050: PAGE <= 12'd296;
            12'd2051: PAGE <= 12'd818;
            12'd2052: PAGE <= 12'd1340;
            12'd2053: PAGE <= 12'd4095;
            12'd2054: PAGE <= 12'd4095;
            12'd2055: PAGE <= 12'd4095;
            12'd2056: PAGE <= 12'd4095;
            12'd2057: PAGE <= 12'd4095;
            12'd2058: PAGE <= 12'd4095;
            12'd2059: PAGE <= 12'd4095;
            12'd2060: PAGE <= 12'd4095;
            12'd2061: PAGE <= 12'd4095;
            12'd2062: PAGE <= 12'd4095;
            12'd2063: PAGE <= 12'd4095;
            12'd2064: PAGE <= 12'd4095;
            12'd2065: PAGE <= 12'd4095;
            12'd2066: PAGE <= 12'd4095;
            12'd2067: PAGE <= 12'd4095;
            12'd2068: PAGE <= 12'd4095;
            12'd2069: PAGE <= 12'd4095;
            12'd2070: PAGE <= 12'd4095;
            12'd2071: PAGE <= 12'd4095;
            12'd2072: PAGE <= 12'd4095;
            12'd2073: PAGE <= 12'd4095;
            12'd2074: PAGE <= 12'd4095;
            12'd2075: PAGE <= 12'd4095;
            12'd2076: PAGE <= 12'd4095;
            12'd2077: PAGE <= 12'd4095;
            12'd2078: PAGE <= 12'd4095;
            12'd2079: PAGE <= 12'd4095;
            12'd2080: PAGE <= 12'd4095;
            12'd2081: PAGE <= 12'd4095;
            12'd2082: PAGE <= 12'd4095;
            12'd2083: PAGE <= 12'd4095;
            12'd2084: PAGE <= 12'd4095;
            12'd2085: PAGE <= 12'd4095;
            12'd2086: PAGE <= 12'd4095;
            12'd2087: PAGE <= 12'd4095;
            12'd2088: PAGE <= 12'd4095;
            12'd2089: PAGE <= 12'd4095;
            12'd2090: PAGE <= 12'd4095;
            12'd2091: PAGE <= 12'd4095;
            12'd2092: PAGE <= 12'd4095;
            12'd2093: PAGE <= 12'd4095;
            12'd2094: PAGE <= 12'd4095;
            12'd2095: PAGE <= 12'd4095;
            12'd2096: PAGE <= 12'd4095;
            12'd2097: PAGE <= 12'd4095;
            12'd2098: PAGE <= 12'd4095;
            12'd2099: PAGE <= 12'd4095;
            12'd2100: PAGE <= 12'd4095;
            12'd2101: PAGE <= 12'd4095;
            12'd2102: PAGE <= 12'd4095;
            12'd2103: PAGE <= 12'd4095;
            12'd2104: PAGE <= 12'd4095;
            12'd2105: PAGE <= 12'd4095;
            12'd2106: PAGE <= 12'd4095;
            12'd2107: PAGE <= 12'd4095;
            12'd2108: PAGE <= 12'd4095;
            12'd2109: PAGE <= 12'd4095;
            12'd2110: PAGE <= 12'd4095;
            12'd2111: PAGE <= 12'd4095;
            12'd2112: PAGE <= 12'd4095;
            12'd2113: PAGE <= 12'd4095;
            12'd2114: PAGE <= 12'd4095;
            12'd2115: PAGE <= 12'd4095;
            12'd2116: PAGE <= 12'd4095;
            12'd2117: PAGE <= 12'd4095;
            12'd2118: PAGE <= 12'd4095;
            12'd2119: PAGE <= 12'd4095;
            12'd2120: PAGE <= 12'd4095;
            12'd2121: PAGE <= 12'd4095;
            12'd2122: PAGE <= 12'd4095;
            12'd2123: PAGE <= 12'd4095;
            12'd2124: PAGE <= 12'd4095;
            12'd2125: PAGE <= 12'd4095;
            12'd2126: PAGE <= 12'd4095;
            12'd2127: PAGE <= 12'd4095;
            12'd2128: PAGE <= 12'd4095;
            12'd2129: PAGE <= 12'd4095;
            12'd2130: PAGE <= 12'd4095;
            12'd2131: PAGE <= 12'd4095;
            12'd2132: PAGE <= 12'd4095;
            12'd2133: PAGE <= 12'd4095;
            12'd2134: PAGE <= 12'd4095;
            12'd2135: PAGE <= 12'd4095;
            12'd2136: PAGE <= 12'd4095;
            12'd2137: PAGE <= 12'd4095;
            12'd2138: PAGE <= 12'd4095;
            12'd2139: PAGE <= 12'd4095;
            12'd2140: PAGE <= 12'd4095;
            12'd2141: PAGE <= 12'd4095;
            12'd2142: PAGE <= 12'd4095;
            12'd2143: PAGE <= 12'd4095;
            12'd2144: PAGE <= 12'd4095;
            12'd2145: PAGE <= 12'd4095;
            12'd2146: PAGE <= 12'd4095;
            12'd2147: PAGE <= 12'd4095;
            12'd2148: PAGE <= 12'd4095;
            12'd2149: PAGE <= 12'd4095;
            12'd2150: PAGE <= 12'd4095;
            12'd2151: PAGE <= 12'd4095;
            12'd2152: PAGE <= 12'd4095;
            12'd2153: PAGE <= 12'd4095;
            12'd2154: PAGE <= 12'd4095;
            12'd2155: PAGE <= 12'd4095;
            12'd2156: PAGE <= 12'd4095;
            12'd2157: PAGE <= 12'd4095;
            12'd2158: PAGE <= 12'd4095;
            12'd2159: PAGE <= 12'd4095;
            12'd2160: PAGE <= 12'd4095;
            12'd2161: PAGE <= 12'd4095;
            12'd2162: PAGE <= 12'd4095;
            12'd2163: PAGE <= 12'd4095;
            12'd2164: PAGE <= 12'd4095;
            12'd2165: PAGE <= 12'd4095;
            12'd2166: PAGE <= 12'd4095;
            12'd2167: PAGE <= 12'd4095;
            12'd2168: PAGE <= 12'd4095;
            12'd2169: PAGE <= 12'd4095;
            12'd2170: PAGE <= 12'd4095;
            12'd2171: PAGE <= 12'd4095;
            12'd2172: PAGE <= 12'd4095;
            12'd2173: PAGE <= 12'd4095;
            12'd2174: PAGE <= 12'd4095;
            12'd2175: PAGE <= 12'd4095;
            12'd2176: PAGE <= 12'd4095;
            12'd2177: PAGE <= 12'd4095;
            12'd2178: PAGE <= 12'd4095;
            12'd2179: PAGE <= 12'd4095;
            12'd2180: PAGE <= 12'd4095;
            12'd2181: PAGE <= 12'd4095;
            12'd2182: PAGE <= 12'd4095;
            12'd2183: PAGE <= 12'd4095;
            12'd2184: PAGE <= 12'd4095;
            12'd2185: PAGE <= 12'd4095;
            12'd2186: PAGE <= 12'd4095;
            12'd2187: PAGE <= 12'd4095;
            12'd2188: PAGE <= 12'd4095;
            12'd2189: PAGE <= 12'd4095;
            12'd2190: PAGE <= 12'd4095;
            12'd2191: PAGE <= 12'd4095;
            12'd2192: PAGE <= 12'd4095;
            12'd2193: PAGE <= 12'd4095;
            12'd2194: PAGE <= 12'd4095;
            12'd2195: PAGE <= 12'd4095;
            12'd2196: PAGE <= 12'd4095;
            12'd2197: PAGE <= 12'd4095;
            12'd2198: PAGE <= 12'd4095;
            12'd2199: PAGE <= 12'd4095;
            12'd2200: PAGE <= 12'd4095;
            12'd2201: PAGE <= 12'd4095;
            12'd2202: PAGE <= 12'd4095;
            12'd2203: PAGE <= 12'd4095;
            12'd2204: PAGE <= 12'd4095;
            12'd2205: PAGE <= 12'd4095;
            12'd2206: PAGE <= 12'd4095;
            12'd2207: PAGE <= 12'd4095;
            12'd2208: PAGE <= 12'd4095;
            12'd2209: PAGE <= 12'd4095;
            12'd2210: PAGE <= 12'd4095;
            12'd2211: PAGE <= 12'd4095;
            12'd2212: PAGE <= 12'd4095;
            12'd2213: PAGE <= 12'd4095;
            12'd2214: PAGE <= 12'd4095;
            12'd2215: PAGE <= 12'd4095;
            12'd2216: PAGE <= 12'd4095;
            12'd2217: PAGE <= 12'd4095;
            12'd2218: PAGE <= 12'd4095;
            12'd2219: PAGE <= 12'd4095;
            12'd2220: PAGE <= 12'd4095;
            12'd2221: PAGE <= 12'd4095;
            12'd2222: PAGE <= 12'd4095;
            12'd2223: PAGE <= 12'd4095;
            12'd2224: PAGE <= 12'd4095;
            12'd2225: PAGE <= 12'd4095;
            12'd2226: PAGE <= 12'd4095;
            12'd2227: PAGE <= 12'd4095;
            12'd2228: PAGE <= 12'd4095;
            12'd2229: PAGE <= 12'd4095;
            12'd2230: PAGE <= 12'd4095;
            12'd2231: PAGE <= 12'd4095;
            12'd2232: PAGE <= 12'd4095;
            12'd2233: PAGE <= 12'd4095;
            12'd2234: PAGE <= 12'd4095;
            12'd2235: PAGE <= 12'd4095;
            12'd2236: PAGE <= 12'd4095;
            12'd2237: PAGE <= 12'd4095;
            12'd2238: PAGE <= 12'd4095;
            12'd2239: PAGE <= 12'd4095;
            12'd2240: PAGE <= 12'd4095;
            12'd2241: PAGE <= 12'd4095;
            12'd2242: PAGE <= 12'd4095;
            12'd2243: PAGE <= 12'd4095;
            12'd2244: PAGE <= 12'd4095;
            12'd2245: PAGE <= 12'd4095;
            12'd2246: PAGE <= 12'd4095;
            12'd2247: PAGE <= 12'd4095;
            12'd2248: PAGE <= 12'd4095;
            12'd2249: PAGE <= 12'd4095;
            12'd2250: PAGE <= 12'd4095;
            12'd2251: PAGE <= 12'd4095;
            12'd2252: PAGE <= 12'd4095;
            12'd2253: PAGE <= 12'd4095;
            12'd2254: PAGE <= 12'd4095;
            12'd2255: PAGE <= 12'd4095;
            12'd2256: PAGE <= 12'd4095;
            12'd2257: PAGE <= 12'd4095;
            12'd2258: PAGE <= 12'd4095;
            12'd2259: PAGE <= 12'd4095;
            12'd2260: PAGE <= 12'd4095;
            12'd2261: PAGE <= 12'd4095;
            12'd2262: PAGE <= 12'd4095;
            12'd2263: PAGE <= 12'd4095;
            12'd2264: PAGE <= 12'd4095;
            12'd2265: PAGE <= 12'd4095;
            12'd2266: PAGE <= 12'd4095;
            12'd2267: PAGE <= 12'd4095;
            12'd2268: PAGE <= 12'd4095;
            12'd2269: PAGE <= 12'd4095;
            12'd2270: PAGE <= 12'd4095;
            12'd2271: PAGE <= 12'd4095;
            12'd2272: PAGE <= 12'd4095;
            12'd2273: PAGE <= 12'd4095;
            12'd2274: PAGE <= 12'd4095;
            12'd2275: PAGE <= 12'd4095;
            12'd2276: PAGE <= 12'd4095;
            12'd2277: PAGE <= 12'd4095;
            12'd2278: PAGE <= 12'd4095;
            12'd2279: PAGE <= 12'd4095;
            12'd2280: PAGE <= 12'd4095;
            12'd2281: PAGE <= 12'd4095;
            12'd2282: PAGE <= 12'd4095;
            12'd2283: PAGE <= 12'd4095;
            12'd2284: PAGE <= 12'd4095;
            12'd2285: PAGE <= 12'd4095;
            12'd2286: PAGE <= 12'd4095;
            12'd2287: PAGE <= 12'd4095;
            12'd2288: PAGE <= 12'd4095;
            12'd2289: PAGE <= 12'd4095;
            12'd2290: PAGE <= 12'd4095;
            12'd2291: PAGE <= 12'd4095;
            12'd2292: PAGE <= 12'd4095;
            12'd2293: PAGE <= 12'd4095;
            12'd2294: PAGE <= 12'd4095;
            12'd2295: PAGE <= 12'd4095;
            12'd2296: PAGE <= 12'd4095;
            12'd2297: PAGE <= 12'd4095;
            12'd2298: PAGE <= 12'd4095;
            12'd2299: PAGE <= 12'd4095;
            12'd2300: PAGE <= 12'd4095;
            12'd2301: PAGE <= 12'd4095;
            12'd2302: PAGE <= 12'd4095;
            12'd2303: PAGE <= 12'd4095;
            12'd2304: PAGE <= 12'd4095;
            12'd2305: PAGE <= 12'd4095;
            12'd2306: PAGE <= 12'd4095;
            12'd2307: PAGE <= 12'd4095;
            12'd2308: PAGE <= 12'd4095;
            12'd2309: PAGE <= 12'd4095;
            12'd2310: PAGE <= 12'd4095;
            12'd2311: PAGE <= 12'd4095;
            12'd2312: PAGE <= 12'd4095;
            12'd2313: PAGE <= 12'd4095;
            12'd2314: PAGE <= 12'd4095;
            12'd2315: PAGE <= 12'd4095;
            12'd2316: PAGE <= 12'd4095;
            12'd2317: PAGE <= 12'd4095;
            12'd2318: PAGE <= 12'd4095;
            12'd2319: PAGE <= 12'd4095;
            12'd2320: PAGE <= 12'd4095;
            12'd2321: PAGE <= 12'd4095;
            12'd2322: PAGE <= 12'd4095;
            12'd2323: PAGE <= 12'd4095;
            12'd2324: PAGE <= 12'd4095;
            12'd2325: PAGE <= 12'd4095;
            12'd2326: PAGE <= 12'd4095;
            12'd2327: PAGE <= 12'd4095;
            12'd2328: PAGE <= 12'd4095;
            12'd2329: PAGE <= 12'd4095;
            12'd2330: PAGE <= 12'd4095;
            12'd2331: PAGE <= 12'd4095;
            12'd2332: PAGE <= 12'd4095;
            12'd2333: PAGE <= 12'd4095;
            12'd2334: PAGE <= 12'd4095;
            12'd2335: PAGE <= 12'd4095;
            12'd2336: PAGE <= 12'd4095;
            12'd2337: PAGE <= 12'd4095;
            12'd2338: PAGE <= 12'd4095;
            12'd2339: PAGE <= 12'd4095;
            12'd2340: PAGE <= 12'd4095;
            12'd2341: PAGE <= 12'd4095;
            12'd2342: PAGE <= 12'd4095;
            12'd2343: PAGE <= 12'd4095;
            12'd2344: PAGE <= 12'd4095;
            12'd2345: PAGE <= 12'd4095;
            12'd2346: PAGE <= 12'd4095;
            12'd2347: PAGE <= 12'd4095;
            12'd2348: PAGE <= 12'd4095;
            12'd2349: PAGE <= 12'd4095;
            12'd2350: PAGE <= 12'd4095;
            12'd2351: PAGE <= 12'd4095;
            12'd2352: PAGE <= 12'd4095;
            12'd2353: PAGE <= 12'd4095;
            12'd2354: PAGE <= 12'd4095;
            12'd2355: PAGE <= 12'd4095;
            12'd2356: PAGE <= 12'd4095;
            12'd2357: PAGE <= 12'd4095;
            12'd2358: PAGE <= 12'd4095;
            12'd2359: PAGE <= 12'd4095;
            12'd2360: PAGE <= 12'd4095;
            12'd2361: PAGE <= 12'd4095;
            12'd2362: PAGE <= 12'd4095;
            12'd2363: PAGE <= 12'd4095;
            12'd2364: PAGE <= 12'd4095;
            12'd2365: PAGE <= 12'd4095;
            12'd2366: PAGE <= 12'd4095;
            12'd2367: PAGE <= 12'd4095;
            12'd2368: PAGE <= 12'd4095;
            12'd2369: PAGE <= 12'd4095;
            12'd2370: PAGE <= 12'd4095;
            12'd2371: PAGE <= 12'd4095;
            12'd2372: PAGE <= 12'd4095;
            12'd2373: PAGE <= 12'd4095;
            12'd2374: PAGE <= 12'd4095;
            12'd2375: PAGE <= 12'd4095;
            12'd2376: PAGE <= 12'd4095;
            12'd2377: PAGE <= 12'd4095;
            12'd2378: PAGE <= 12'd4095;
            12'd2379: PAGE <= 12'd4095;
            12'd2380: PAGE <= 12'd4095;
            12'd2381: PAGE <= 12'd4095;
            12'd2382: PAGE <= 12'd4095;
            12'd2383: PAGE <= 12'd4095;
            12'd2384: PAGE <= 12'd4095;
            12'd2385: PAGE <= 12'd4095;
            12'd2386: PAGE <= 12'd4095;
            12'd2387: PAGE <= 12'd4095;
            12'd2388: PAGE <= 12'd4095;
            12'd2389: PAGE <= 12'd4095;
            12'd2390: PAGE <= 12'd4095;
            12'd2391: PAGE <= 12'd4095;
            12'd2392: PAGE <= 12'd4095;
            12'd2393: PAGE <= 12'd4095;
            12'd2394: PAGE <= 12'd4095;
            12'd2395: PAGE <= 12'd4095;
            12'd2396: PAGE <= 12'd4095;
            12'd2397: PAGE <= 12'd4095;
            12'd2398: PAGE <= 12'd4095;
            12'd2399: PAGE <= 12'd4095;
            12'd2400: PAGE <= 12'd4095;
            12'd2401: PAGE <= 12'd4095;
            12'd2402: PAGE <= 12'd4095;
            12'd2403: PAGE <= 12'd4095;
            12'd2404: PAGE <= 12'd4095;
            12'd2405: PAGE <= 12'd4095;
            12'd2406: PAGE <= 12'd4095;
            12'd2407: PAGE <= 12'd4095;
            12'd2408: PAGE <= 12'd4095;
            12'd2409: PAGE <= 12'd4095;
            12'd2410: PAGE <= 12'd4095;
            12'd2411: PAGE <= 12'd4095;
            12'd2412: PAGE <= 12'd4095;
            12'd2413: PAGE <= 12'd4095;
            12'd2414: PAGE <= 12'd4095;
            12'd2415: PAGE <= 12'd4095;
            12'd2416: PAGE <= 12'd4095;
            12'd2417: PAGE <= 12'd4095;
            12'd2418: PAGE <= 12'd4095;
            12'd2419: PAGE <= 12'd4095;
            12'd2420: PAGE <= 12'd4095;
            12'd2421: PAGE <= 12'd4095;
            12'd2422: PAGE <= 12'd4095;
            12'd2423: PAGE <= 12'd4095;
            12'd2424: PAGE <= 12'd4095;
            12'd2425: PAGE <= 12'd4095;
            12'd2426: PAGE <= 12'd4095;
            12'd2427: PAGE <= 12'd4095;
            12'd2428: PAGE <= 12'd4095;
            12'd2429: PAGE <= 12'd4095;
            12'd2430: PAGE <= 12'd4095;
            12'd2431: PAGE <= 12'd4095;
            12'd2432: PAGE <= 12'd4095;
            12'd2433: PAGE <= 12'd4095;
            12'd2434: PAGE <= 12'd4095;
            12'd2435: PAGE <= 12'd4095;
            12'd2436: PAGE <= 12'd4095;
            12'd2437: PAGE <= 12'd4095;
            12'd2438: PAGE <= 12'd4095;
            12'd2439: PAGE <= 12'd4095;
            12'd2440: PAGE <= 12'd4095;
            12'd2441: PAGE <= 12'd4095;
            12'd2442: PAGE <= 12'd4095;
            12'd2443: PAGE <= 12'd4095;
            12'd2444: PAGE <= 12'd4095;
            12'd2445: PAGE <= 12'd4095;
            12'd2446: PAGE <= 12'd4095;
            12'd2447: PAGE <= 12'd4095;
            12'd2448: PAGE <= 12'd4095;
            12'd2449: PAGE <= 12'd4095;
            12'd2450: PAGE <= 12'd4095;
            12'd2451: PAGE <= 12'd4095;
            12'd2452: PAGE <= 12'd4095;
            12'd2453: PAGE <= 12'd4095;
            12'd2454: PAGE <= 12'd4095;
            12'd2455: PAGE <= 12'd4095;
            12'd2456: PAGE <= 12'd4095;
            12'd2457: PAGE <= 12'd4095;
            12'd2458: PAGE <= 12'd4095;
            12'd2459: PAGE <= 12'd4095;
            12'd2460: PAGE <= 12'd4095;
            12'd2461: PAGE <= 12'd4095;
            12'd2462: PAGE <= 12'd4095;
            12'd2463: PAGE <= 12'd4095;
            12'd2464: PAGE <= 12'd4095;
            12'd2465: PAGE <= 12'd4095;
            12'd2466: PAGE <= 12'd4095;
            12'd2467: PAGE <= 12'd4095;
            12'd2468: PAGE <= 12'd4095;
            12'd2469: PAGE <= 12'd4095;
            12'd2470: PAGE <= 12'd4095;
            12'd2471: PAGE <= 12'd4095;
            12'd2472: PAGE <= 12'd4095;
            12'd2473: PAGE <= 12'd4095;
            12'd2474: PAGE <= 12'd4095;
            12'd2475: PAGE <= 12'd4095;
            12'd2476: PAGE <= 12'd4095;
            12'd2477: PAGE <= 12'd4095;
            12'd2478: PAGE <= 12'd4095;
            12'd2479: PAGE <= 12'd4095;
            12'd2480: PAGE <= 12'd4095;
            12'd2481: PAGE <= 12'd4095;
            12'd2482: PAGE <= 12'd4095;
            12'd2483: PAGE <= 12'd4095;
            12'd2484: PAGE <= 12'd4095;
            12'd2485: PAGE <= 12'd4095;
            12'd2486: PAGE <= 12'd4095;
            12'd2487: PAGE <= 12'd4095;
            12'd2488: PAGE <= 12'd4095;
            12'd2489: PAGE <= 12'd4095;
            12'd2490: PAGE <= 12'd4095;
            12'd2491: PAGE <= 12'd4095;
            12'd2492: PAGE <= 12'd4095;
            12'd2493: PAGE <= 12'd4095;
            12'd2494: PAGE <= 12'd4095;
            12'd2495: PAGE <= 12'd4095;
            12'd2496: PAGE <= 12'd4095;
            12'd2497: PAGE <= 12'd4095;
            12'd2498: PAGE <= 12'd4095;
            12'd2499: PAGE <= 12'd4095;
            12'd2500: PAGE <= 12'd4095;
            12'd2501: PAGE <= 12'd4095;
            12'd2502: PAGE <= 12'd4095;
            12'd2503: PAGE <= 12'd4095;
            12'd2504: PAGE <= 12'd4095;
            12'd2505: PAGE <= 12'd4095;
            12'd2506: PAGE <= 12'd4095;
            12'd2507: PAGE <= 12'd4095;
            12'd2508: PAGE <= 12'd4095;
            12'd2509: PAGE <= 12'd4095;
            12'd2510: PAGE <= 12'd4095;
            12'd2511: PAGE <= 12'd4095;
            12'd2512: PAGE <= 12'd4095;
            12'd2513: PAGE <= 12'd4095;
            12'd2514: PAGE <= 12'd4095;
            12'd2515: PAGE <= 12'd4095;
            12'd2516: PAGE <= 12'd4095;
            12'd2517: PAGE <= 12'd4095;
            12'd2518: PAGE <= 12'd4095;
            12'd2519: PAGE <= 12'd4095;
            12'd2520: PAGE <= 12'd4095;
            12'd2521: PAGE <= 12'd4095;
            12'd2522: PAGE <= 12'd4095;
            12'd2523: PAGE <= 12'd4095;
            12'd2524: PAGE <= 12'd4095;
            12'd2525: PAGE <= 12'd4095;
            12'd2526: PAGE <= 12'd4095;
            12'd2527: PAGE <= 12'd4095;
            12'd2528: PAGE <= 12'd4095;
            12'd2529: PAGE <= 12'd4095;
            12'd2530: PAGE <= 12'd4095;
            12'd2531: PAGE <= 12'd4095;
            12'd2532: PAGE <= 12'd4095;
            12'd2533: PAGE <= 12'd4095;
            12'd2534: PAGE <= 12'd4095;
            12'd2535: PAGE <= 12'd4095;
            12'd2536: PAGE <= 12'd4095;
            12'd2537: PAGE <= 12'd4095;
            12'd2538: PAGE <= 12'd4095;
            12'd2539: PAGE <= 12'd4095;
            12'd2540: PAGE <= 12'd4095;
            12'd2541: PAGE <= 12'd4095;
            12'd2542: PAGE <= 12'd4095;
            12'd2543: PAGE <= 12'd4095;
            12'd2544: PAGE <= 12'd4095;
            12'd2545: PAGE <= 12'd4095;
            12'd2546: PAGE <= 12'd4095;
            12'd2547: PAGE <= 12'd4095;
            12'd2548: PAGE <= 12'd4095;
            12'd2549: PAGE <= 12'd4095;
            12'd2550: PAGE <= 12'd4095;
            12'd2551: PAGE <= 12'd4095;
            12'd2552: PAGE <= 12'd4095;
            12'd2553: PAGE <= 12'd4095;
            12'd2554: PAGE <= 12'd4095;
            12'd2555: PAGE <= 12'd4095;
            12'd2556: PAGE <= 12'd4095;
            12'd2557: PAGE <= 12'd4095;
            12'd2558: PAGE <= 12'd4095;
            12'd2559: PAGE <= 12'd4095;
            12'd2560: PAGE <= 12'd4095;
            12'd2561: PAGE <= 12'd4095;
            12'd2562: PAGE <= 12'd4095;
            12'd2563: PAGE <= 12'd4095;
            12'd2564: PAGE <= 12'd4095;
            12'd2565: PAGE <= 12'd4095;
            12'd2566: PAGE <= 12'd4095;
            12'd2567: PAGE <= 12'd4095;
            12'd2568: PAGE <= 12'd4095;
            12'd2569: PAGE <= 12'd4095;
            12'd2570: PAGE <= 12'd4095;
            12'd2571: PAGE <= 12'd4095;
            12'd2572: PAGE <= 12'd4095;
            12'd2573: PAGE <= 12'd4095;
            12'd2574: PAGE <= 12'd4095;
            12'd2575: PAGE <= 12'd4095;
            12'd2576: PAGE <= 12'd4095;
            12'd2577: PAGE <= 12'd4095;
            12'd2578: PAGE <= 12'd4095;
            12'd2579: PAGE <= 12'd4095;
            12'd2580: PAGE <= 12'd4095;
            12'd2581: PAGE <= 12'd4095;
            12'd2582: PAGE <= 12'd4095;
            12'd2583: PAGE <= 12'd4095;
            12'd2584: PAGE <= 12'd4095;
            12'd2585: PAGE <= 12'd4095;
            12'd2586: PAGE <= 12'd4095;
            12'd2587: PAGE <= 12'd4095;
            12'd2588: PAGE <= 12'd4095;
            12'd2589: PAGE <= 12'd4095;
            12'd2590: PAGE <= 12'd4095;
            12'd2591: PAGE <= 12'd4095;
            12'd2592: PAGE <= 12'd4095;
            12'd2593: PAGE <= 12'd4095;
            12'd2594: PAGE <= 12'd4095;
            12'd2595: PAGE <= 12'd4095;
            12'd2596: PAGE <= 12'd4095;
            12'd2597: PAGE <= 12'd4095;
            12'd2598: PAGE <= 12'd4095;
            12'd2599: PAGE <= 12'd4095;
            12'd2600: PAGE <= 12'd4095;
            12'd2601: PAGE <= 12'd4095;
            12'd2602: PAGE <= 12'd4095;
            12'd2603: PAGE <= 12'd4095;
            12'd2604: PAGE <= 12'd4095;
            12'd2605: PAGE <= 12'd4095;
            12'd2606: PAGE <= 12'd4095;
            12'd2607: PAGE <= 12'd4095;
            12'd2608: PAGE <= 12'd4095;
            12'd2609: PAGE <= 12'd4095;
            12'd2610: PAGE <= 12'd4095;
            12'd2611: PAGE <= 12'd4095;
            12'd2612: PAGE <= 12'd4095;
            12'd2613: PAGE <= 12'd4095;
            12'd2614: PAGE <= 12'd4095;
            12'd2615: PAGE <= 12'd4095;
            12'd2616: PAGE <= 12'd4095;
            12'd2617: PAGE <= 12'd4095;
            12'd2618: PAGE <= 12'd4095;
            12'd2619: PAGE <= 12'd4095;
            12'd2620: PAGE <= 12'd4095;
            12'd2621: PAGE <= 12'd4095;
            12'd2622: PAGE <= 12'd4095;
            12'd2623: PAGE <= 12'd4095;
            12'd2624: PAGE <= 12'd4095;
            12'd2625: PAGE <= 12'd4095;
            12'd2626: PAGE <= 12'd4095;
            12'd2627: PAGE <= 12'd4095;
            12'd2628: PAGE <= 12'd4095;
            12'd2629: PAGE <= 12'd4095;
            12'd2630: PAGE <= 12'd4095;
            12'd2631: PAGE <= 12'd4095;
            12'd2632: PAGE <= 12'd4095;
            12'd2633: PAGE <= 12'd4095;
            12'd2634: PAGE <= 12'd4095;
            12'd2635: PAGE <= 12'd4095;
            12'd2636: PAGE <= 12'd4095;
            12'd2637: PAGE <= 12'd4095;
            12'd2638: PAGE <= 12'd4095;
            12'd2639: PAGE <= 12'd4095;
            12'd2640: PAGE <= 12'd4095;
            12'd2641: PAGE <= 12'd4095;
            12'd2642: PAGE <= 12'd4095;
            12'd2643: PAGE <= 12'd4095;
            12'd2644: PAGE <= 12'd4095;
            12'd2645: PAGE <= 12'd4095;
            12'd2646: PAGE <= 12'd4095;
            12'd2647: PAGE <= 12'd4095;
            12'd2648: PAGE <= 12'd4095;
            12'd2649: PAGE <= 12'd4095;
            12'd2650: PAGE <= 12'd4095;
            12'd2651: PAGE <= 12'd4095;
            12'd2652: PAGE <= 12'd4095;
            12'd2653: PAGE <= 12'd4095;
            12'd2654: PAGE <= 12'd4095;
            12'd2655: PAGE <= 12'd4095;
            12'd2656: PAGE <= 12'd4095;
            12'd2657: PAGE <= 12'd4095;
            12'd2658: PAGE <= 12'd4095;
            12'd2659: PAGE <= 12'd4095;
            12'd2660: PAGE <= 12'd4095;
            12'd2661: PAGE <= 12'd4095;
            12'd2662: PAGE <= 12'd4095;
            12'd2663: PAGE <= 12'd4095;
            12'd2664: PAGE <= 12'd4095;
            12'd2665: PAGE <= 12'd4095;
            12'd2666: PAGE <= 12'd4095;
            12'd2667: PAGE <= 12'd4095;
            12'd2668: PAGE <= 12'd4095;
            12'd2669: PAGE <= 12'd4095;
            12'd2670: PAGE <= 12'd4095;
            12'd2671: PAGE <= 12'd4095;
            12'd2672: PAGE <= 12'd4095;
            12'd2673: PAGE <= 12'd4095;
            12'd2674: PAGE <= 12'd4095;
            12'd2675: PAGE <= 12'd4095;
            12'd2676: PAGE <= 12'd4095;
            12'd2677: PAGE <= 12'd4095;
            12'd2678: PAGE <= 12'd4095;
            12'd2679: PAGE <= 12'd4095;
            12'd2680: PAGE <= 12'd4095;
            12'd2681: PAGE <= 12'd4095;
            12'd2682: PAGE <= 12'd4095;
            12'd2683: PAGE <= 12'd4095;
            12'd2684: PAGE <= 12'd4095;
            12'd2685: PAGE <= 12'd4095;
            12'd2686: PAGE <= 12'd4095;
            12'd2687: PAGE <= 12'd4095;
            12'd2688: PAGE <= 12'd4095;
            12'd2689: PAGE <= 12'd4095;
            12'd2690: PAGE <= 12'd4095;
            12'd2691: PAGE <= 12'd4095;
            12'd2692: PAGE <= 12'd4095;
            12'd2693: PAGE <= 12'd4095;
            12'd2694: PAGE <= 12'd4095;
            12'd2695: PAGE <= 12'd4095;
            12'd2696: PAGE <= 12'd4095;
            12'd2697: PAGE <= 12'd4095;
            12'd2698: PAGE <= 12'd4095;
            12'd2699: PAGE <= 12'd4095;
            12'd2700: PAGE <= 12'd4095;
            12'd2701: PAGE <= 12'd4095;
            12'd2702: PAGE <= 12'd4095;
            12'd2703: PAGE <= 12'd4095;
            12'd2704: PAGE <= 12'd4095;
            12'd2705: PAGE <= 12'd4095;
            12'd2706: PAGE <= 12'd4095;
            12'd2707: PAGE <= 12'd4095;
            12'd2708: PAGE <= 12'd4095;
            12'd2709: PAGE <= 12'd4095;
            12'd2710: PAGE <= 12'd4095;
            12'd2711: PAGE <= 12'd4095;
            12'd2712: PAGE <= 12'd4095;
            12'd2713: PAGE <= 12'd4095;
            12'd2714: PAGE <= 12'd4095;
            12'd2715: PAGE <= 12'd4095;
            12'd2716: PAGE <= 12'd4095;
            12'd2717: PAGE <= 12'd4095;
            12'd2718: PAGE <= 12'd4095;
            12'd2719: PAGE <= 12'd4095;
            12'd2720: PAGE <= 12'd4095;
            12'd2721: PAGE <= 12'd4095;
            12'd2722: PAGE <= 12'd4095;
            12'd2723: PAGE <= 12'd4095;
            12'd2724: PAGE <= 12'd4095;
            12'd2725: PAGE <= 12'd4095;
            12'd2726: PAGE <= 12'd4095;
            12'd2727: PAGE <= 12'd4095;
            12'd2728: PAGE <= 12'd4095;
            12'd2729: PAGE <= 12'd4095;
            12'd2730: PAGE <= 12'd4095;
            12'd2731: PAGE <= 12'd4095;
            12'd2732: PAGE <= 12'd4095;
            12'd2733: PAGE <= 12'd4095;
            12'd2734: PAGE <= 12'd4095;
            12'd2735: PAGE <= 12'd4095;
            12'd2736: PAGE <= 12'd4095;
            12'd2737: PAGE <= 12'd4095;
            12'd2738: PAGE <= 12'd4095;
            12'd2739: PAGE <= 12'd4095;
            12'd2740: PAGE <= 12'd4095;
            12'd2741: PAGE <= 12'd4095;
            12'd2742: PAGE <= 12'd4095;
            12'd2743: PAGE <= 12'd4095;
            12'd2744: PAGE <= 12'd4095;
            12'd2745: PAGE <= 12'd4095;
            12'd2746: PAGE <= 12'd4095;
            12'd2747: PAGE <= 12'd4095;
            12'd2748: PAGE <= 12'd4095;
            12'd2749: PAGE <= 12'd4095;
            12'd2750: PAGE <= 12'd4095;
            12'd2751: PAGE <= 12'd4095;
            12'd2752: PAGE <= 12'd4095;
            12'd2753: PAGE <= 12'd4095;
            12'd2754: PAGE <= 12'd4095;
            12'd2755: PAGE <= 12'd4095;
            12'd2756: PAGE <= 12'd4095;
            12'd2757: PAGE <= 12'd4095;
            12'd2758: PAGE <= 12'd4095;
            12'd2759: PAGE <= 12'd4095;
            12'd2760: PAGE <= 12'd4095;
            12'd2761: PAGE <= 12'd4095;
            12'd2762: PAGE <= 12'd4095;
            12'd2763: PAGE <= 12'd4095;
            12'd2764: PAGE <= 12'd4095;
            12'd2765: PAGE <= 12'd4095;
            12'd2766: PAGE <= 12'd4095;
            12'd2767: PAGE <= 12'd4095;
            12'd2768: PAGE <= 12'd4095;
            12'd2769: PAGE <= 12'd4095;
            12'd2770: PAGE <= 12'd4095;
            12'd2771: PAGE <= 12'd4095;
            12'd2772: PAGE <= 12'd4095;
            12'd2773: PAGE <= 12'd4095;
            12'd2774: PAGE <= 12'd4095;
            12'd2775: PAGE <= 12'd4095;
            12'd2776: PAGE <= 12'd4095;
            12'd2777: PAGE <= 12'd4095;
            12'd2778: PAGE <= 12'd4095;
            12'd2779: PAGE <= 12'd4095;
            12'd2780: PAGE <= 12'd4095;
            12'd2781: PAGE <= 12'd4095;
            12'd2782: PAGE <= 12'd4095;
            12'd2783: PAGE <= 12'd4095;
            12'd2784: PAGE <= 12'd4095;
            12'd2785: PAGE <= 12'd4095;
            12'd2786: PAGE <= 12'd4095;
            12'd2787: PAGE <= 12'd4095;
            12'd2788: PAGE <= 12'd4095;
            12'd2789: PAGE <= 12'd4095;
            12'd2790: PAGE <= 12'd4095;
            12'd2791: PAGE <= 12'd4095;
            12'd2792: PAGE <= 12'd4095;
            12'd2793: PAGE <= 12'd4095;
            12'd2794: PAGE <= 12'd4095;
            12'd2795: PAGE <= 12'd4095;
            12'd2796: PAGE <= 12'd4095;
            12'd2797: PAGE <= 12'd4095;
            12'd2798: PAGE <= 12'd4095;
            12'd2799: PAGE <= 12'd4095;
            12'd2800: PAGE <= 12'd4095;
            12'd2801: PAGE <= 12'd4095;
            12'd2802: PAGE <= 12'd4095;
            12'd2803: PAGE <= 12'd4095;
            12'd2804: PAGE <= 12'd4095;
            12'd2805: PAGE <= 12'd4095;
            12'd2806: PAGE <= 12'd4095;
            12'd2807: PAGE <= 12'd4095;
            12'd2808: PAGE <= 12'd4095;
            12'd2809: PAGE <= 12'd4095;
            12'd2810: PAGE <= 12'd4095;
            12'd2811: PAGE <= 12'd4095;
            12'd2812: PAGE <= 12'd4095;
            12'd2813: PAGE <= 12'd4095;
            12'd2814: PAGE <= 12'd4095;
            12'd2815: PAGE <= 12'd4095;
            12'd2816: PAGE <= 12'd4095;
            12'd2817: PAGE <= 12'd4095;
            12'd2818: PAGE <= 12'd4095;
            12'd2819: PAGE <= 12'd4095;
            12'd2820: PAGE <= 12'd4095;
            12'd2821: PAGE <= 12'd4095;
            12'd2822: PAGE <= 12'd4095;
            12'd2823: PAGE <= 12'd4095;
            12'd2824: PAGE <= 12'd4095;
            12'd2825: PAGE <= 12'd4095;
            12'd2826: PAGE <= 12'd4095;
            12'd2827: PAGE <= 12'd4095;
            12'd2828: PAGE <= 12'd4095;
            12'd2829: PAGE <= 12'd4095;
            12'd2830: PAGE <= 12'd4095;
            12'd2831: PAGE <= 12'd4095;
            12'd2832: PAGE <= 12'd4095;
            12'd2833: PAGE <= 12'd4095;
            12'd2834: PAGE <= 12'd4095;
            12'd2835: PAGE <= 12'd4095;
            12'd2836: PAGE <= 12'd4095;
            12'd2837: PAGE <= 12'd4095;
            12'd2838: PAGE <= 12'd4095;
            12'd2839: PAGE <= 12'd4095;
            12'd2840: PAGE <= 12'd4095;
            12'd2841: PAGE <= 12'd4095;
            12'd2842: PAGE <= 12'd4095;
            12'd2843: PAGE <= 12'd4095;
            12'd2844: PAGE <= 12'd4095;
            12'd2845: PAGE <= 12'd4095;
            12'd2846: PAGE <= 12'd4095;
            12'd2847: PAGE <= 12'd4095;
            12'd2848: PAGE <= 12'd4095;
            12'd2849: PAGE <= 12'd4095;
            12'd2850: PAGE <= 12'd4095;
            12'd2851: PAGE <= 12'd4095;
            12'd2852: PAGE <= 12'd4095;
            12'd2853: PAGE <= 12'd4095;
            12'd2854: PAGE <= 12'd4095;
            12'd2855: PAGE <= 12'd4095;
            12'd2856: PAGE <= 12'd4095;
            12'd2857: PAGE <= 12'd4095;
            12'd2858: PAGE <= 12'd4095;
            12'd2859: PAGE <= 12'd4095;
            12'd2860: PAGE <= 12'd4095;
            12'd2861: PAGE <= 12'd4095;
            12'd2862: PAGE <= 12'd4095;
            12'd2863: PAGE <= 12'd4095;
            12'd2864: PAGE <= 12'd4095;
            12'd2865: PAGE <= 12'd4095;
            12'd2866: PAGE <= 12'd4095;
            12'd2867: PAGE <= 12'd4095;
            12'd2868: PAGE <= 12'd4095;
            12'd2869: PAGE <= 12'd4095;
            12'd2870: PAGE <= 12'd4095;
            12'd2871: PAGE <= 12'd4095;
            12'd2872: PAGE <= 12'd4095;
            12'd2873: PAGE <= 12'd4095;
            12'd2874: PAGE <= 12'd4095;
            12'd2875: PAGE <= 12'd4095;
            12'd2876: PAGE <= 12'd4095;
            12'd2877: PAGE <= 12'd4095;
            12'd2878: PAGE <= 12'd4095;
            12'd2879: PAGE <= 12'd4095;
            12'd2880: PAGE <= 12'd4095;
            12'd2881: PAGE <= 12'd4095;
            12'd2882: PAGE <= 12'd4095;
            12'd2883: PAGE <= 12'd4095;
            12'd2884: PAGE <= 12'd4095;
            12'd2885: PAGE <= 12'd4095;
            12'd2886: PAGE <= 12'd4095;
            12'd2887: PAGE <= 12'd4095;
            12'd2888: PAGE <= 12'd4095;
            12'd2889: PAGE <= 12'd4095;
            12'd2890: PAGE <= 12'd4095;
            12'd2891: PAGE <= 12'd4095;
            12'd2892: PAGE <= 12'd4095;
            12'd2893: PAGE <= 12'd4095;
            12'd2894: PAGE <= 12'd4095;
            12'd2895: PAGE <= 12'd4095;
            12'd2896: PAGE <= 12'd4095;
            12'd2897: PAGE <= 12'd4095;
            12'd2898: PAGE <= 12'd4095;
            12'd2899: PAGE <= 12'd4095;
            12'd2900: PAGE <= 12'd4095;
            12'd2901: PAGE <= 12'd4095;
            12'd2902: PAGE <= 12'd4095;
            12'd2903: PAGE <= 12'd4095;
            12'd2904: PAGE <= 12'd4095;
            12'd2905: PAGE <= 12'd4095;
            12'd2906: PAGE <= 12'd4095;
            12'd2907: PAGE <= 12'd4095;
            12'd2908: PAGE <= 12'd4095;
            12'd2909: PAGE <= 12'd4095;
            12'd2910: PAGE <= 12'd4095;
            12'd2911: PAGE <= 12'd4095;
            12'd2912: PAGE <= 12'd4095;
            12'd2913: PAGE <= 12'd4095;
            12'd2914: PAGE <= 12'd4095;
            12'd2915: PAGE <= 12'd4095;
            12'd2916: PAGE <= 12'd4095;
            12'd2917: PAGE <= 12'd4095;
            12'd2918: PAGE <= 12'd4095;
            12'd2919: PAGE <= 12'd4095;
            12'd2920: PAGE <= 12'd4095;
            12'd2921: PAGE <= 12'd4095;
            12'd2922: PAGE <= 12'd4095;
            12'd2923: PAGE <= 12'd4095;
            12'd2924: PAGE <= 12'd4095;
            12'd2925: PAGE <= 12'd4095;
            12'd2926: PAGE <= 12'd4095;
            12'd2927: PAGE <= 12'd4095;
            12'd2928: PAGE <= 12'd4095;
            12'd2929: PAGE <= 12'd4095;
            12'd2930: PAGE <= 12'd4095;
            12'd2931: PAGE <= 12'd4095;
            12'd2932: PAGE <= 12'd4095;
            12'd2933: PAGE <= 12'd4095;
            12'd2934: PAGE <= 12'd4095;
            12'd2935: PAGE <= 12'd4095;
            12'd2936: PAGE <= 12'd4095;
            12'd2937: PAGE <= 12'd4095;
            12'd2938: PAGE <= 12'd4095;
            12'd2939: PAGE <= 12'd4095;
            12'd2940: PAGE <= 12'd4095;
            12'd2941: PAGE <= 12'd4095;
            12'd2942: PAGE <= 12'd4095;
            12'd2943: PAGE <= 12'd4095;
            12'd2944: PAGE <= 12'd4095;
            12'd2945: PAGE <= 12'd4095;
            12'd2946: PAGE <= 12'd4095;
            12'd2947: PAGE <= 12'd4095;
            12'd2948: PAGE <= 12'd4095;
            12'd2949: PAGE <= 12'd4095;
            12'd2950: PAGE <= 12'd4095;
            12'd2951: PAGE <= 12'd4095;
            12'd2952: PAGE <= 12'd4095;
            12'd2953: PAGE <= 12'd4095;
            12'd2954: PAGE <= 12'd4095;
            12'd2955: PAGE <= 12'd4095;
            12'd2956: PAGE <= 12'd4095;
            12'd2957: PAGE <= 12'd4095;
            12'd2958: PAGE <= 12'd4095;
            12'd2959: PAGE <= 12'd4095;
            12'd2960: PAGE <= 12'd4095;
            12'd2961: PAGE <= 12'd4095;
            12'd2962: PAGE <= 12'd4095;
            12'd2963: PAGE <= 12'd4095;
            12'd2964: PAGE <= 12'd4095;
            12'd2965: PAGE <= 12'd4095;
            12'd2966: PAGE <= 12'd4095;
            12'd2967: PAGE <= 12'd4095;
            12'd2968: PAGE <= 12'd4095;
            12'd2969: PAGE <= 12'd4095;
            12'd2970: PAGE <= 12'd4095;
            12'd2971: PAGE <= 12'd4095;
            12'd2972: PAGE <= 12'd4095;
            12'd2973: PAGE <= 12'd4095;
            12'd2974: PAGE <= 12'd4095;
            12'd2975: PAGE <= 12'd4095;
            12'd2976: PAGE <= 12'd4095;
            12'd2977: PAGE <= 12'd4095;
            12'd2978: PAGE <= 12'd4095;
            12'd2979: PAGE <= 12'd4095;
            12'd2980: PAGE <= 12'd4095;
            12'd2981: PAGE <= 12'd4095;
            12'd2982: PAGE <= 12'd4095;
            12'd2983: PAGE <= 12'd4095;
            12'd2984: PAGE <= 12'd4095;
            12'd2985: PAGE <= 12'd4095;
            12'd2986: PAGE <= 12'd4095;
            12'd2987: PAGE <= 12'd4095;
            12'd2988: PAGE <= 12'd4095;
            12'd2989: PAGE <= 12'd4095;
            12'd2990: PAGE <= 12'd4095;
            12'd2991: PAGE <= 12'd4095;
            12'd2992: PAGE <= 12'd4095;
            12'd2993: PAGE <= 12'd4095;
            12'd2994: PAGE <= 12'd4095;
            12'd2995: PAGE <= 12'd4095;
            12'd2996: PAGE <= 12'd4095;
            12'd2997: PAGE <= 12'd4095;
            12'd2998: PAGE <= 12'd4095;
            12'd2999: PAGE <= 12'd4095;
            12'd3000: PAGE <= 12'd4095;
            12'd3001: PAGE <= 12'd4095;
            12'd3002: PAGE <= 12'd4095;
            12'd3003: PAGE <= 12'd4095;
            12'd3004: PAGE <= 12'd4095;
            12'd3005: PAGE <= 12'd4095;
            12'd3006: PAGE <= 12'd4095;
            12'd3007: PAGE <= 12'd4095;
            12'd3008: PAGE <= 12'd4095;
            12'd3009: PAGE <= 12'd4095;
            12'd3010: PAGE <= 12'd4095;
            12'd3011: PAGE <= 12'd4095;
            12'd3012: PAGE <= 12'd4095;
            12'd3013: PAGE <= 12'd4095;
            12'd3014: PAGE <= 12'd4095;
            12'd3015: PAGE <= 12'd4095;
            12'd3016: PAGE <= 12'd4095;
            12'd3017: PAGE <= 12'd4095;
            12'd3018: PAGE <= 12'd4095;
            12'd3019: PAGE <= 12'd4095;
            12'd3020: PAGE <= 12'd4095;
            12'd3021: PAGE <= 12'd4095;
            12'd3022: PAGE <= 12'd4095;
            12'd3023: PAGE <= 12'd4095;
            12'd3024: PAGE <= 12'd4095;
            12'd3025: PAGE <= 12'd4095;
            12'd3026: PAGE <= 12'd4095;
            12'd3027: PAGE <= 12'd4095;
            12'd3028: PAGE <= 12'd4095;
            12'd3029: PAGE <= 12'd4095;
            12'd3030: PAGE <= 12'd4095;
            12'd3031: PAGE <= 12'd4095;
            12'd3032: PAGE <= 12'd4095;
            12'd3033: PAGE <= 12'd4095;
            12'd3034: PAGE <= 12'd4095;
            12'd3035: PAGE <= 12'd4095;
            12'd3036: PAGE <= 12'd4095;
            12'd3037: PAGE <= 12'd4095;
            12'd3038: PAGE <= 12'd4095;
            12'd3039: PAGE <= 12'd4095;
            12'd3040: PAGE <= 12'd4095;
            12'd3041: PAGE <= 12'd4095;
            12'd3042: PAGE <= 12'd4095;
            12'd3043: PAGE <= 12'd4095;
            12'd3044: PAGE <= 12'd4095;
            12'd3045: PAGE <= 12'd4095;
            12'd3046: PAGE <= 12'd4095;
            12'd3047: PAGE <= 12'd4095;
            12'd3048: PAGE <= 12'd4095;
            12'd3049: PAGE <= 12'd4095;
            12'd3050: PAGE <= 12'd4095;
            12'd3051: PAGE <= 12'd4095;
            12'd3052: PAGE <= 12'd4095;
            12'd3053: PAGE <= 12'd4095;
            12'd3054: PAGE <= 12'd4095;
            12'd3055: PAGE <= 12'd4095;
            12'd3056: PAGE <= 12'd4095;
            12'd3057: PAGE <= 12'd4095;
            12'd3058: PAGE <= 12'd4095;
            12'd3059: PAGE <= 12'd4095;
            12'd3060: PAGE <= 12'd4095;
            12'd3061: PAGE <= 12'd4095;
            12'd3062: PAGE <= 12'd4095;
            12'd3063: PAGE <= 12'd4095;
            12'd3064: PAGE <= 12'd4095;
            12'd3065: PAGE <= 12'd4095;
            12'd3066: PAGE <= 12'd4095;
            12'd3067: PAGE <= 12'd4095;
            12'd3068: PAGE <= 12'd4095;
            12'd3069: PAGE <= 12'd4095;
            12'd3070: PAGE <= 12'd4095;
            12'd3071: PAGE <= 12'd4095;
            12'd3072: PAGE <= 12'd4095;
            12'd3073: PAGE <= 12'd4095;
            12'd3074: PAGE <= 12'd4095;
            12'd3075: PAGE <= 12'd4095;
            12'd3076: PAGE <= 12'd4095;
            12'd3077: PAGE <= 12'd4095;
            12'd3078: PAGE <= 12'd4095;
            12'd3079: PAGE <= 12'd4095;
            12'd3080: PAGE <= 12'd4095;
            12'd3081: PAGE <= 12'd4095;
            12'd3082: PAGE <= 12'd4095;
            12'd3083: PAGE <= 12'd4095;
            12'd3084: PAGE <= 12'd4095;
            12'd3085: PAGE <= 12'd4095;
            12'd3086: PAGE <= 12'd4095;
            12'd3087: PAGE <= 12'd4095;
            12'd3088: PAGE <= 12'd4095;
            12'd3089: PAGE <= 12'd4095;
            12'd3090: PAGE <= 12'd4095;
            12'd3091: PAGE <= 12'd4095;
            12'd3092: PAGE <= 12'd4095;
            12'd3093: PAGE <= 12'd4095;
            12'd3094: PAGE <= 12'd4095;
            12'd3095: PAGE <= 12'd4095;
            12'd3096: PAGE <= 12'd4095;
            12'd3097: PAGE <= 12'd4095;
            12'd3098: PAGE <= 12'd4095;
            12'd3099: PAGE <= 12'd4095;
            12'd3100: PAGE <= 12'd4095;
            12'd3101: PAGE <= 12'd4095;
            12'd3102: PAGE <= 12'd4095;
            12'd3103: PAGE <= 12'd4095;
            12'd3104: PAGE <= 12'd4095;
            12'd3105: PAGE <= 12'd4095;
            12'd3106: PAGE <= 12'd4095;
            12'd3107: PAGE <= 12'd4095;
            12'd3108: PAGE <= 12'd4095;
            12'd3109: PAGE <= 12'd4095;
            12'd3110: PAGE <= 12'd4095;
            12'd3111: PAGE <= 12'd4095;
            12'd3112: PAGE <= 12'd4095;
            12'd3113: PAGE <= 12'd4095;
            12'd3114: PAGE <= 12'd4095;
            12'd3115: PAGE <= 12'd4095;
            12'd3116: PAGE <= 12'd4095;
            12'd3117: PAGE <= 12'd4095;
            12'd3118: PAGE <= 12'd4095;
            12'd3119: PAGE <= 12'd4095;
            12'd3120: PAGE <= 12'd4095;
            12'd3121: PAGE <= 12'd4095;
            12'd3122: PAGE <= 12'd4095;
            12'd3123: PAGE <= 12'd4095;
            12'd3124: PAGE <= 12'd4095;
            12'd3125: PAGE <= 12'd4095;
            12'd3126: PAGE <= 12'd4095;
            12'd3127: PAGE <= 12'd4095;
            12'd3128: PAGE <= 12'd4095;
            12'd3129: PAGE <= 12'd4095;
            12'd3130: PAGE <= 12'd4095;
            12'd3131: PAGE <= 12'd4095;
            12'd3132: PAGE <= 12'd4095;
            12'd3133: PAGE <= 12'd4095;
            12'd3134: PAGE <= 12'd4095;
            12'd3135: PAGE <= 12'd4095;
            12'd3136: PAGE <= 12'd4095;
            12'd3137: PAGE <= 12'd4095;
            12'd3138: PAGE <= 12'd4095;
            12'd3139: PAGE <= 12'd4095;
            12'd3140: PAGE <= 12'd4095;
            12'd3141: PAGE <= 12'd4095;
            12'd3142: PAGE <= 12'd4095;
            12'd3143: PAGE <= 12'd4095;
            12'd3144: PAGE <= 12'd4095;
            12'd3145: PAGE <= 12'd4095;
            12'd3146: PAGE <= 12'd4095;
            12'd3147: PAGE <= 12'd4095;
            12'd3148: PAGE <= 12'd4095;
            12'd3149: PAGE <= 12'd4095;
            12'd3150: PAGE <= 12'd4095;
            12'd3151: PAGE <= 12'd4095;
            12'd3152: PAGE <= 12'd4095;
            12'd3153: PAGE <= 12'd4095;
            12'd3154: PAGE <= 12'd4095;
            12'd3155: PAGE <= 12'd4095;
            12'd3156: PAGE <= 12'd4095;
            12'd3157: PAGE <= 12'd4095;
            12'd3158: PAGE <= 12'd4095;
            12'd3159: PAGE <= 12'd4095;
            12'd3160: PAGE <= 12'd4095;
            12'd3161: PAGE <= 12'd4095;
            12'd3162: PAGE <= 12'd4095;
            12'd3163: PAGE <= 12'd4095;
            12'd3164: PAGE <= 12'd4095;
            12'd3165: PAGE <= 12'd4095;
            12'd3166: PAGE <= 12'd4095;
            12'd3167: PAGE <= 12'd4095;
            12'd3168: PAGE <= 12'd4095;
            12'd3169: PAGE <= 12'd4095;
            12'd3170: PAGE <= 12'd4095;
            12'd3171: PAGE <= 12'd4095;
            12'd3172: PAGE <= 12'd4095;
            12'd3173: PAGE <= 12'd4095;
            12'd3174: PAGE <= 12'd4095;
            12'd3175: PAGE <= 12'd4095;
            12'd3176: PAGE <= 12'd4095;
            12'd3177: PAGE <= 12'd4095;
            12'd3178: PAGE <= 12'd4095;
            12'd3179: PAGE <= 12'd4095;
            12'd3180: PAGE <= 12'd4095;
            12'd3181: PAGE <= 12'd4095;
            12'd3182: PAGE <= 12'd4095;
            12'd3183: PAGE <= 12'd4095;
            12'd3184: PAGE <= 12'd4095;
            12'd3185: PAGE <= 12'd4095;
            12'd3186: PAGE <= 12'd4095;
            12'd3187: PAGE <= 12'd4095;
            12'd3188: PAGE <= 12'd4095;
            12'd3189: PAGE <= 12'd4095;
            12'd3190: PAGE <= 12'd4095;
            12'd3191: PAGE <= 12'd4095;
            12'd3192: PAGE <= 12'd4095;
            12'd3193: PAGE <= 12'd4095;
            12'd3194: PAGE <= 12'd4095;
            12'd3195: PAGE <= 12'd4095;
            12'd3196: PAGE <= 12'd4095;
            12'd3197: PAGE <= 12'd4095;
            12'd3198: PAGE <= 12'd4095;
            12'd3199: PAGE <= 12'd4095;
            12'd3200: PAGE <= 12'd4095;
            12'd3201: PAGE <= 12'd4095;
            12'd3202: PAGE <= 12'd4095;
            12'd3203: PAGE <= 12'd4095;
            12'd3204: PAGE <= 12'd4095;
            12'd3205: PAGE <= 12'd4095;
            12'd3206: PAGE <= 12'd4095;
            12'd3207: PAGE <= 12'd4095;
            12'd3208: PAGE <= 12'd4095;
            12'd3209: PAGE <= 12'd4095;
            12'd3210: PAGE <= 12'd4095;
            12'd3211: PAGE <= 12'd4095;
            12'd3212: PAGE <= 12'd4095;
            12'd3213: PAGE <= 12'd4095;
            12'd3214: PAGE <= 12'd4095;
            12'd3215: PAGE <= 12'd4095;
            12'd3216: PAGE <= 12'd4095;
            12'd3217: PAGE <= 12'd4095;
            12'd3218: PAGE <= 12'd4095;
            12'd3219: PAGE <= 12'd4095;
            12'd3220: PAGE <= 12'd4095;
            12'd3221: PAGE <= 12'd4095;
            12'd3222: PAGE <= 12'd4095;
            12'd3223: PAGE <= 12'd4095;
            12'd3224: PAGE <= 12'd4095;
            12'd3225: PAGE <= 12'd4095;
            12'd3226: PAGE <= 12'd4095;
            12'd3227: PAGE <= 12'd4095;
            12'd3228: PAGE <= 12'd4095;
            12'd3229: PAGE <= 12'd4095;
            12'd3230: PAGE <= 12'd4095;
            12'd3231: PAGE <= 12'd4095;
            12'd3232: PAGE <= 12'd4095;
            12'd3233: PAGE <= 12'd4095;
            12'd3234: PAGE <= 12'd4095;
            12'd3235: PAGE <= 12'd4095;
            12'd3236: PAGE <= 12'd4095;
            12'd3237: PAGE <= 12'd4095;
            12'd3238: PAGE <= 12'd4095;
            12'd3239: PAGE <= 12'd4095;
            12'd3240: PAGE <= 12'd4095;
            12'd3241: PAGE <= 12'd4095;
            12'd3242: PAGE <= 12'd4095;
            12'd3243: PAGE <= 12'd4095;
            12'd3244: PAGE <= 12'd4095;
            12'd3245: PAGE <= 12'd4095;
            12'd3246: PAGE <= 12'd4095;
            12'd3247: PAGE <= 12'd4095;
            12'd3248: PAGE <= 12'd4095;
            12'd3249: PAGE <= 12'd4095;
            12'd3250: PAGE <= 12'd4095;
            12'd3251: PAGE <= 12'd4095;
            12'd3252: PAGE <= 12'd4095;
            12'd3253: PAGE <= 12'd4095;
            12'd3254: PAGE <= 12'd4095;
            12'd3255: PAGE <= 12'd4095;
            12'd3256: PAGE <= 12'd4095;
            12'd3257: PAGE <= 12'd4095;
            12'd3258: PAGE <= 12'd4095;
            12'd3259: PAGE <= 12'd4095;
            12'd3260: PAGE <= 12'd4095;
            12'd3261: PAGE <= 12'd4095;
            12'd3262: PAGE <= 12'd4095;
            12'd3263: PAGE <= 12'd4095;
            12'd3264: PAGE <= 12'd4095;
            12'd3265: PAGE <= 12'd4095;
            12'd3266: PAGE <= 12'd4095;
            12'd3267: PAGE <= 12'd4095;
            12'd3268: PAGE <= 12'd4095;
            12'd3269: PAGE <= 12'd4095;
            12'd3270: PAGE <= 12'd4095;
            12'd3271: PAGE <= 12'd4095;
            12'd3272: PAGE <= 12'd4095;
            12'd3273: PAGE <= 12'd4095;
            12'd3274: PAGE <= 12'd4095;
            12'd3275: PAGE <= 12'd4095;
            12'd3276: PAGE <= 12'd4095;
            12'd3277: PAGE <= 12'd4095;
            12'd3278: PAGE <= 12'd4095;
            12'd3279: PAGE <= 12'd4095;
            12'd3280: PAGE <= 12'd4095;
            12'd3281: PAGE <= 12'd4095;
            12'd3282: PAGE <= 12'd4095;
            12'd3283: PAGE <= 12'd4095;
            12'd3284: PAGE <= 12'd4095;
            12'd3285: PAGE <= 12'd4095;
            12'd3286: PAGE <= 12'd4095;
            12'd3287: PAGE <= 12'd4095;
            12'd3288: PAGE <= 12'd4095;
            12'd3289: PAGE <= 12'd4095;
            12'd3290: PAGE <= 12'd4095;
            12'd3291: PAGE <= 12'd4095;
            12'd3292: PAGE <= 12'd4095;
            12'd3293: PAGE <= 12'd4095;
            12'd3294: PAGE <= 12'd4095;
            12'd3295: PAGE <= 12'd4095;
            12'd3296: PAGE <= 12'd4095;
            12'd3297: PAGE <= 12'd4095;
            12'd3298: PAGE <= 12'd4095;
            12'd3299: PAGE <= 12'd4095;
            12'd3300: PAGE <= 12'd4095;
            12'd3301: PAGE <= 12'd4095;
            12'd3302: PAGE <= 12'd4095;
            12'd3303: PAGE <= 12'd4095;
            12'd3304: PAGE <= 12'd4095;
            12'd3305: PAGE <= 12'd4095;
            12'd3306: PAGE <= 12'd4095;
            12'd3307: PAGE <= 12'd4095;
            12'd3308: PAGE <= 12'd4095;
            12'd3309: PAGE <= 12'd4095;
            12'd3310: PAGE <= 12'd4095;
            12'd3311: PAGE <= 12'd4095;
            12'd3312: PAGE <= 12'd4095;
            12'd3313: PAGE <= 12'd4095;
            12'd3314: PAGE <= 12'd4095;
            12'd3315: PAGE <= 12'd4095;
            12'd3316: PAGE <= 12'd4095;
            12'd3317: PAGE <= 12'd4095;
            12'd3318: PAGE <= 12'd4095;
            12'd3319: PAGE <= 12'd4095;
            12'd3320: PAGE <= 12'd4095;
            12'd3321: PAGE <= 12'd4095;
            12'd3322: PAGE <= 12'd4095;
            12'd3323: PAGE <= 12'd4095;
            12'd3324: PAGE <= 12'd4095;
            12'd3325: PAGE <= 12'd4095;
            12'd3326: PAGE <= 12'd4095;
            12'd3327: PAGE <= 12'd4095;
            12'd3328: PAGE <= 12'd4095;
            12'd3329: PAGE <= 12'd4095;
            12'd3330: PAGE <= 12'd4095;
            12'd3331: PAGE <= 12'd4095;
            12'd3332: PAGE <= 12'd4095;
            12'd3333: PAGE <= 12'd4095;
            12'd3334: PAGE <= 12'd4095;
            12'd3335: PAGE <= 12'd4095;
            12'd3336: PAGE <= 12'd4095;
            12'd3337: PAGE <= 12'd4095;
            12'd3338: PAGE <= 12'd4095;
            12'd3339: PAGE <= 12'd4095;
            12'd3340: PAGE <= 12'd4095;
            12'd3341: PAGE <= 12'd4095;
            12'd3342: PAGE <= 12'd4095;
            12'd3343: PAGE <= 12'd4095;
            12'd3344: PAGE <= 12'd4095;
            12'd3345: PAGE <= 12'd4095;
            12'd3346: PAGE <= 12'd4095;
            12'd3347: PAGE <= 12'd4095;
            12'd3348: PAGE <= 12'd4095;
            12'd3349: PAGE <= 12'd4095;
            12'd3350: PAGE <= 12'd4095;
            12'd3351: PAGE <= 12'd4095;
            12'd3352: PAGE <= 12'd4095;
            12'd3353: PAGE <= 12'd4095;
            12'd3354: PAGE <= 12'd4095;
            12'd3355: PAGE <= 12'd4095;
            12'd3356: PAGE <= 12'd4095;
            12'd3357: PAGE <= 12'd4095;
            12'd3358: PAGE <= 12'd4095;
            12'd3359: PAGE <= 12'd4095;
            12'd3360: PAGE <= 12'd4095;
            12'd3361: PAGE <= 12'd4095;
            12'd3362: PAGE <= 12'd4095;
            12'd3363: PAGE <= 12'd4095;
            12'd3364: PAGE <= 12'd4095;
            12'd3365: PAGE <= 12'd4095;
            12'd3366: PAGE <= 12'd4095;
            12'd3367: PAGE <= 12'd4095;
            12'd3368: PAGE <= 12'd4095;
            12'd3369: PAGE <= 12'd4095;
            12'd3370: PAGE <= 12'd4095;
            12'd3371: PAGE <= 12'd4095;
            12'd3372: PAGE <= 12'd4095;
            12'd3373: PAGE <= 12'd4095;
            12'd3374: PAGE <= 12'd4095;
            12'd3375: PAGE <= 12'd4095;
            12'd3376: PAGE <= 12'd4095;
            12'd3377: PAGE <= 12'd4095;
            12'd3378: PAGE <= 12'd4095;
            12'd3379: PAGE <= 12'd4095;
            12'd3380: PAGE <= 12'd4095;
            12'd3381: PAGE <= 12'd4095;
            12'd3382: PAGE <= 12'd4095;
            12'd3383: PAGE <= 12'd4095;
            12'd3384: PAGE <= 12'd4095;
            12'd3385: PAGE <= 12'd4095;
            12'd3386: PAGE <= 12'd4095;
            12'd3387: PAGE <= 12'd4095;
            12'd3388: PAGE <= 12'd4095;
            12'd3389: PAGE <= 12'd4095;
            12'd3390: PAGE <= 12'd4095;
            12'd3391: PAGE <= 12'd4095;
            12'd3392: PAGE <= 12'd4095;
            12'd3393: PAGE <= 12'd4095;
            12'd3394: PAGE <= 12'd4095;
            12'd3395: PAGE <= 12'd4095;
            12'd3396: PAGE <= 12'd4095;
            12'd3397: PAGE <= 12'd4095;
            12'd3398: PAGE <= 12'd4095;
            12'd3399: PAGE <= 12'd4095;
            12'd3400: PAGE <= 12'd4095;
            12'd3401: PAGE <= 12'd4095;
            12'd3402: PAGE <= 12'd4095;
            12'd3403: PAGE <= 12'd4095;
            12'd3404: PAGE <= 12'd4095;
            12'd3405: PAGE <= 12'd4095;
            12'd3406: PAGE <= 12'd4095;
            12'd3407: PAGE <= 12'd4095;
            12'd3408: PAGE <= 12'd4095;
            12'd3409: PAGE <= 12'd4095;
            12'd3410: PAGE <= 12'd4095;
            12'd3411: PAGE <= 12'd4095;
            12'd3412: PAGE <= 12'd4095;
            12'd3413: PAGE <= 12'd4095;
            12'd3414: PAGE <= 12'd4095;
            12'd3415: PAGE <= 12'd4095;
            12'd3416: PAGE <= 12'd4095;
            12'd3417: PAGE <= 12'd4095;
            12'd3418: PAGE <= 12'd4095;
            12'd3419: PAGE <= 12'd4095;
            12'd3420: PAGE <= 12'd4095;
            12'd3421: PAGE <= 12'd4095;
            12'd3422: PAGE <= 12'd4095;
            12'd3423: PAGE <= 12'd4095;
            12'd3424: PAGE <= 12'd4095;
            12'd3425: PAGE <= 12'd4095;
            12'd3426: PAGE <= 12'd4095;
            12'd3427: PAGE <= 12'd4095;
            12'd3428: PAGE <= 12'd4095;
            12'd3429: PAGE <= 12'd4095;
            12'd3430: PAGE <= 12'd4095;
            12'd3431: PAGE <= 12'd4095;
            12'd3432: PAGE <= 12'd4095;
            12'd3433: PAGE <= 12'd4095;
            12'd3434: PAGE <= 12'd4095;
            12'd3435: PAGE <= 12'd4095;
            12'd3436: PAGE <= 12'd4095;
            12'd3437: PAGE <= 12'd4095;
            12'd3438: PAGE <= 12'd4095;
            12'd3439: PAGE <= 12'd4095;
            12'd3440: PAGE <= 12'd4095;
            12'd3441: PAGE <= 12'd4095;
            12'd3442: PAGE <= 12'd4095;
            12'd3443: PAGE <= 12'd4095;
            12'd3444: PAGE <= 12'd4095;
            12'd3445: PAGE <= 12'd4095;
            12'd3446: PAGE <= 12'd4095;
            12'd3447: PAGE <= 12'd4095;
            12'd3448: PAGE <= 12'd4095;
            12'd3449: PAGE <= 12'd4095;
            12'd3450: PAGE <= 12'd4095;
            12'd3451: PAGE <= 12'd4095;
            12'd3452: PAGE <= 12'd4095;
            12'd3453: PAGE <= 12'd4095;
            12'd3454: PAGE <= 12'd4095;
            12'd3455: PAGE <= 12'd4095;
            12'd3456: PAGE <= 12'd4095;
            12'd3457: PAGE <= 12'd4095;
            12'd3458: PAGE <= 12'd4095;
            12'd3459: PAGE <= 12'd4095;
            12'd3460: PAGE <= 12'd4095;
            12'd3461: PAGE <= 12'd4095;
            12'd3462: PAGE <= 12'd4095;
            12'd3463: PAGE <= 12'd4095;
            12'd3464: PAGE <= 12'd4095;
            12'd3465: PAGE <= 12'd4095;
            12'd3466: PAGE <= 12'd4095;
            12'd3467: PAGE <= 12'd4095;
            12'd3468: PAGE <= 12'd4095;
            12'd3469: PAGE <= 12'd4095;
            12'd3470: PAGE <= 12'd4095;
            12'd3471: PAGE <= 12'd4095;
            12'd3472: PAGE <= 12'd4095;
            12'd3473: PAGE <= 12'd4095;
            12'd3474: PAGE <= 12'd4095;
            12'd3475: PAGE <= 12'd4095;
            12'd3476: PAGE <= 12'd4095;
            12'd3477: PAGE <= 12'd4095;
            12'd3478: PAGE <= 12'd4095;
            12'd3479: PAGE <= 12'd4095;
            12'd3480: PAGE <= 12'd4095;
            12'd3481: PAGE <= 12'd4095;
            12'd3482: PAGE <= 12'd4095;
            12'd3483: PAGE <= 12'd4095;
            12'd3484: PAGE <= 12'd4095;
            12'd3485: PAGE <= 12'd4095;
            12'd3486: PAGE <= 12'd4095;
            12'd3487: PAGE <= 12'd4095;
            12'd3488: PAGE <= 12'd4095;
            12'd3489: PAGE <= 12'd4095;
            12'd3490: PAGE <= 12'd4095;
            12'd3491: PAGE <= 12'd4095;
            12'd3492: PAGE <= 12'd4095;
            12'd3493: PAGE <= 12'd4095;
            12'd3494: PAGE <= 12'd4095;
            12'd3495: PAGE <= 12'd4095;
            12'd3496: PAGE <= 12'd4095;
            12'd3497: PAGE <= 12'd4095;
            12'd3498: PAGE <= 12'd4095;
            12'd3499: PAGE <= 12'd4095;
            12'd3500: PAGE <= 12'd4095;
            12'd3501: PAGE <= 12'd4095;
            12'd3502: PAGE <= 12'd4095;
            12'd3503: PAGE <= 12'd4095;
            12'd3504: PAGE <= 12'd4095;
            12'd3505: PAGE <= 12'd4095;
            12'd3506: PAGE <= 12'd4095;
            12'd3507: PAGE <= 12'd4095;
            12'd3508: PAGE <= 12'd4095;
            12'd3509: PAGE <= 12'd4095;
            12'd3510: PAGE <= 12'd4095;
            12'd3511: PAGE <= 12'd4095;
            12'd3512: PAGE <= 12'd4095;
            12'd3513: PAGE <= 12'd4095;
            12'd3514: PAGE <= 12'd4095;
            12'd3515: PAGE <= 12'd4095;
            12'd3516: PAGE <= 12'd4095;
            12'd3517: PAGE <= 12'd4095;
            12'd3518: PAGE <= 12'd4095;
            12'd3519: PAGE <= 12'd4095;
            12'd3520: PAGE <= 12'd4095;
            12'd3521: PAGE <= 12'd4095;
            12'd3522: PAGE <= 12'd4095;
            12'd3523: PAGE <= 12'd4095;
            12'd3524: PAGE <= 12'd4095;
            12'd3525: PAGE <= 12'd4095;
            12'd3526: PAGE <= 12'd4095;
            12'd3527: PAGE <= 12'd4095;
            12'd3528: PAGE <= 12'd4095;
            12'd3529: PAGE <= 12'd4095;
            12'd3530: PAGE <= 12'd4095;
            12'd3531: PAGE <= 12'd4095;
            12'd3532: PAGE <= 12'd4095;
            12'd3533: PAGE <= 12'd4095;
            12'd3534: PAGE <= 12'd4095;
            12'd3535: PAGE <= 12'd4095;
            12'd3536: PAGE <= 12'd4095;
            12'd3537: PAGE <= 12'd4095;
            12'd3538: PAGE <= 12'd4095;
            12'd3539: PAGE <= 12'd4095;
            12'd3540: PAGE <= 12'd4095;
            12'd3541: PAGE <= 12'd4095;
            12'd3542: PAGE <= 12'd4095;
            12'd3543: PAGE <= 12'd4095;
            12'd3544: PAGE <= 12'd4095;
            12'd3545: PAGE <= 12'd4095;
            12'd3546: PAGE <= 12'd4095;
            12'd3547: PAGE <= 12'd4095;
            12'd3548: PAGE <= 12'd4095;
            12'd3549: PAGE <= 12'd4095;
            12'd3550: PAGE <= 12'd4095;
            12'd3551: PAGE <= 12'd4095;
            12'd3552: PAGE <= 12'd4095;
            12'd3553: PAGE <= 12'd4095;
            12'd3554: PAGE <= 12'd4095;
            12'd3555: PAGE <= 12'd4095;
            12'd3556: PAGE <= 12'd4095;
            12'd3557: PAGE <= 12'd4095;
            12'd3558: PAGE <= 12'd4095;
            12'd3559: PAGE <= 12'd4095;
            12'd3560: PAGE <= 12'd4095;
            12'd3561: PAGE <= 12'd4095;
            12'd3562: PAGE <= 12'd4095;
            12'd3563: PAGE <= 12'd4095;
            12'd3564: PAGE <= 12'd4095;
            12'd3565: PAGE <= 12'd4095;
            12'd3566: PAGE <= 12'd4095;
            12'd3567: PAGE <= 12'd4095;
            12'd3568: PAGE <= 12'd4095;
            12'd3569: PAGE <= 12'd4095;
            12'd3570: PAGE <= 12'd4095;
            12'd3571: PAGE <= 12'd4095;
            12'd3572: PAGE <= 12'd4095;
            12'd3573: PAGE <= 12'd4095;
            12'd3574: PAGE <= 12'd4095;
            12'd3575: PAGE <= 12'd4095;
            12'd3576: PAGE <= 12'd4095;
            12'd3577: PAGE <= 12'd4095;
            12'd3578: PAGE <= 12'd4095;
            12'd3579: PAGE <= 12'd4095;
            12'd3580: PAGE <= 12'd4095;
            12'd3581: PAGE <= 12'd4095;
            12'd3582: PAGE <= 12'd4095;
            12'd3583: PAGE <= 12'd4095;
            12'd3584: PAGE <= 12'd4095;
            12'd3585: PAGE <= 12'd4095;
            12'd3586: PAGE <= 12'd4095;
            12'd3587: PAGE <= 12'd4095;
            12'd3588: PAGE <= 12'd4095;
            12'd3589: PAGE <= 12'd4095;
            12'd3590: PAGE <= 12'd4095;
            12'd3591: PAGE <= 12'd4095;
            12'd3592: PAGE <= 12'd4095;
            12'd3593: PAGE <= 12'd4095;
            12'd3594: PAGE <= 12'd4095;
            12'd3595: PAGE <= 12'd4095;
            12'd3596: PAGE <= 12'd4095;
            12'd3597: PAGE <= 12'd4095;
            12'd3598: PAGE <= 12'd4095;
            12'd3599: PAGE <= 12'd4095;
            12'd3600: PAGE <= 12'd4095;
            12'd3601: PAGE <= 12'd4095;
            12'd3602: PAGE <= 12'd4095;
            12'd3603: PAGE <= 12'd4095;
            12'd3604: PAGE <= 12'd4095;
            12'd3605: PAGE <= 12'd4095;
            12'd3606: PAGE <= 12'd4095;
            12'd3607: PAGE <= 12'd4095;
            12'd3608: PAGE <= 12'd4095;
            12'd3609: PAGE <= 12'd4095;
            12'd3610: PAGE <= 12'd4095;
            12'd3611: PAGE <= 12'd4095;
            12'd3612: PAGE <= 12'd4095;
            12'd3613: PAGE <= 12'd4095;
            12'd3614: PAGE <= 12'd4095;
            12'd3615: PAGE <= 12'd4095;
            12'd3616: PAGE <= 12'd4095;
            12'd3617: PAGE <= 12'd4095;
            12'd3618: PAGE <= 12'd4095;
            12'd3619: PAGE <= 12'd4095;
            12'd3620: PAGE <= 12'd4095;
            12'd3621: PAGE <= 12'd4095;
            12'd3622: PAGE <= 12'd4095;
            12'd3623: PAGE <= 12'd4095;
            12'd3624: PAGE <= 12'd4095;
            12'd3625: PAGE <= 12'd4095;
            12'd3626: PAGE <= 12'd4095;
            12'd3627: PAGE <= 12'd4095;
            12'd3628: PAGE <= 12'd4095;
            12'd3629: PAGE <= 12'd4095;
            12'd3630: PAGE <= 12'd4095;
            12'd3631: PAGE <= 12'd4095;
            12'd3632: PAGE <= 12'd4095;
            12'd3633: PAGE <= 12'd4095;
            12'd3634: PAGE <= 12'd4095;
            12'd3635: PAGE <= 12'd4095;
            12'd3636: PAGE <= 12'd4095;
            12'd3637: PAGE <= 12'd4095;
            12'd3638: PAGE <= 12'd4095;
            12'd3639: PAGE <= 12'd4095;
            12'd3640: PAGE <= 12'd4095;
            12'd3641: PAGE <= 12'd4095;
            12'd3642: PAGE <= 12'd4095;
            12'd3643: PAGE <= 12'd4095;
            12'd3644: PAGE <= 12'd4095;
            12'd3645: PAGE <= 12'd4095;
            12'd3646: PAGE <= 12'd4095;
            12'd3647: PAGE <= 12'd4095;
            12'd3648: PAGE <= 12'd4095;
            12'd3649: PAGE <= 12'd4095;
            12'd3650: PAGE <= 12'd4095;
            12'd3651: PAGE <= 12'd4095;
            12'd3652: PAGE <= 12'd4095;
            12'd3653: PAGE <= 12'd4095;
            12'd3654: PAGE <= 12'd4095;
            12'd3655: PAGE <= 12'd4095;
            12'd3656: PAGE <= 12'd4095;
            12'd3657: PAGE <= 12'd4095;
            12'd3658: PAGE <= 12'd4095;
            12'd3659: PAGE <= 12'd4095;
            12'd3660: PAGE <= 12'd4095;
            12'd3661: PAGE <= 12'd4095;
            12'd3662: PAGE <= 12'd4095;
            12'd3663: PAGE <= 12'd4095;
            12'd3664: PAGE <= 12'd4095;
            12'd3665: PAGE <= 12'd4095;
            12'd3666: PAGE <= 12'd4095;
            12'd3667: PAGE <= 12'd4095;
            12'd3668: PAGE <= 12'd4095;
            12'd3669: PAGE <= 12'd4095;
            12'd3670: PAGE <= 12'd4095;
            12'd3671: PAGE <= 12'd4095;
            12'd3672: PAGE <= 12'd4095;
            12'd3673: PAGE <= 12'd4095;
            12'd3674: PAGE <= 12'd4095;
            12'd3675: PAGE <= 12'd4095;
            12'd3676: PAGE <= 12'd4095;
            12'd3677: PAGE <= 12'd4095;
            12'd3678: PAGE <= 12'd4095;
            12'd3679: PAGE <= 12'd4095;
            12'd3680: PAGE <= 12'd4095;
            12'd3681: PAGE <= 12'd4095;
            12'd3682: PAGE <= 12'd4095;
            12'd3683: PAGE <= 12'd4095;
            12'd3684: PAGE <= 12'd4095;
            12'd3685: PAGE <= 12'd4095;
            12'd3686: PAGE <= 12'd4095;
            12'd3687: PAGE <= 12'd4095;
            12'd3688: PAGE <= 12'd4095;
            12'd3689: PAGE <= 12'd4095;
            12'd3690: PAGE <= 12'd4095;
            12'd3691: PAGE <= 12'd4095;
            12'd3692: PAGE <= 12'd4095;
            12'd3693: PAGE <= 12'd4095;
            12'd3694: PAGE <= 12'd4095;
            12'd3695: PAGE <= 12'd4095;
            12'd3696: PAGE <= 12'd4095;
            12'd3697: PAGE <= 12'd4095;
            12'd3698: PAGE <= 12'd4095;
            12'd3699: PAGE <= 12'd4095;
            12'd3700: PAGE <= 12'd4095;
            12'd3701: PAGE <= 12'd4095;
            12'd3702: PAGE <= 12'd4095;
            12'd3703: PAGE <= 12'd4095;
            12'd3704: PAGE <= 12'd4095;
            12'd3705: PAGE <= 12'd4095;
            12'd3706: PAGE <= 12'd4095;
            12'd3707: PAGE <= 12'd4095;
            12'd3708: PAGE <= 12'd4095;
            12'd3709: PAGE <= 12'd4095;
            12'd3710: PAGE <= 12'd4095;
            12'd3711: PAGE <= 12'd4095;
            12'd3712: PAGE <= 12'd4095;
            12'd3713: PAGE <= 12'd4095;
            12'd3714: PAGE <= 12'd4095;
            12'd3715: PAGE <= 12'd4095;
            12'd3716: PAGE <= 12'd4095;
            12'd3717: PAGE <= 12'd4095;
            12'd3718: PAGE <= 12'd4095;
            12'd3719: PAGE <= 12'd4095;
            12'd3720: PAGE <= 12'd4095;
            12'd3721: PAGE <= 12'd4095;
            12'd3722: PAGE <= 12'd4095;
            12'd3723: PAGE <= 12'd4095;
            12'd3724: PAGE <= 12'd4095;
            12'd3725: PAGE <= 12'd4095;
            12'd3726: PAGE <= 12'd4095;
            12'd3727: PAGE <= 12'd4095;
            12'd3728: PAGE <= 12'd4095;
            12'd3729: PAGE <= 12'd4095;
            12'd3730: PAGE <= 12'd4095;
            12'd3731: PAGE <= 12'd4095;
            12'd3732: PAGE <= 12'd4095;
            12'd3733: PAGE <= 12'd4095;
            12'd3734: PAGE <= 12'd4095;
            12'd3735: PAGE <= 12'd4095;
            12'd3736: PAGE <= 12'd4095;
            12'd3737: PAGE <= 12'd4095;
            12'd3738: PAGE <= 12'd4095;
            12'd3739: PAGE <= 12'd4095;
            12'd3740: PAGE <= 12'd4095;
            12'd3741: PAGE <= 12'd4095;
            12'd3742: PAGE <= 12'd4095;
            12'd3743: PAGE <= 12'd4095;
            12'd3744: PAGE <= 12'd4095;
            12'd3745: PAGE <= 12'd4095;
            12'd3746: PAGE <= 12'd4095;
            12'd3747: PAGE <= 12'd4095;
            12'd3748: PAGE <= 12'd4095;
            12'd3749: PAGE <= 12'd4095;
            12'd3750: PAGE <= 12'd4095;
            12'd3751: PAGE <= 12'd4095;
            12'd3752: PAGE <= 12'd4095;
            12'd3753: PAGE <= 12'd4095;
            12'd3754: PAGE <= 12'd4095;
            12'd3755: PAGE <= 12'd4095;
            12'd3756: PAGE <= 12'd4095;
            12'd3757: PAGE <= 12'd4095;
            12'd3758: PAGE <= 12'd4095;
            12'd3759: PAGE <= 12'd4095;
            12'd3760: PAGE <= 12'd4095;
            12'd3761: PAGE <= 12'd4095;
            12'd3762: PAGE <= 12'd4095;
            12'd3763: PAGE <= 12'd4095;
            12'd3764: PAGE <= 12'd4095;
            12'd3765: PAGE <= 12'd4095;
            12'd3766: PAGE <= 12'd4095;
            12'd3767: PAGE <= 12'd4095;
            12'd3768: PAGE <= 12'd4095;
            12'd3769: PAGE <= 12'd4095;
            12'd3770: PAGE <= 12'd4095;
            12'd3771: PAGE <= 12'd4095;
            12'd3772: PAGE <= 12'd4095;
            12'd3773: PAGE <= 12'd4095;
            12'd3774: PAGE <= 12'd4095;
            12'd3775: PAGE <= 12'd4095;
            12'd3776: PAGE <= 12'd4095;
            12'd3777: PAGE <= 12'd4095;
            12'd3778: PAGE <= 12'd4095;
            12'd3779: PAGE <= 12'd4095;
            12'd3780: PAGE <= 12'd4095;
            12'd3781: PAGE <= 12'd4095;
            12'd3782: PAGE <= 12'd4095;
            12'd3783: PAGE <= 12'd4095;
            12'd3784: PAGE <= 12'd4095;
            12'd3785: PAGE <= 12'd4095;
            12'd3786: PAGE <= 12'd4095;
            12'd3787: PAGE <= 12'd4095;
            12'd3788: PAGE <= 12'd4095;
            12'd3789: PAGE <= 12'd4095;
            12'd3790: PAGE <= 12'd4095;
            12'd3791: PAGE <= 12'd4095;
            12'd3792: PAGE <= 12'd4095;
            12'd3793: PAGE <= 12'd4095;
            12'd3794: PAGE <= 12'd4095;
            12'd3795: PAGE <= 12'd4095;
            12'd3796: PAGE <= 12'd4095;
            12'd3797: PAGE <= 12'd4095;
            12'd3798: PAGE <= 12'd4095;
            12'd3799: PAGE <= 12'd4095;
            12'd3800: PAGE <= 12'd4095;
            12'd3801: PAGE <= 12'd4095;
            12'd3802: PAGE <= 12'd4095;
            12'd3803: PAGE <= 12'd4095;
            12'd3804: PAGE <= 12'd4095;
            12'd3805: PAGE <= 12'd4095;
            12'd3806: PAGE <= 12'd4095;
            12'd3807: PAGE <= 12'd4095;
            12'd3808: PAGE <= 12'd4095;
            12'd3809: PAGE <= 12'd4095;
            12'd3810: PAGE <= 12'd4095;
            12'd3811: PAGE <= 12'd4095;
            12'd3812: PAGE <= 12'd4095;
            12'd3813: PAGE <= 12'd4095;
            12'd3814: PAGE <= 12'd4095;
            12'd3815: PAGE <= 12'd4095;
            12'd3816: PAGE <= 12'd4095;
            12'd3817: PAGE <= 12'd4095;
            12'd3818: PAGE <= 12'd4095;
            12'd3819: PAGE <= 12'd4095;
            12'd3820: PAGE <= 12'd4095;
            12'd3821: PAGE <= 12'd4095;
            12'd3822: PAGE <= 12'd4095;
            12'd3823: PAGE <= 12'd4095;
            12'd3824: PAGE <= 12'd4095;
            12'd3825: PAGE <= 12'd4095;
            12'd3826: PAGE <= 12'd4095;
            12'd3827: PAGE <= 12'd4095;
            12'd3828: PAGE <= 12'd4095;
            12'd3829: PAGE <= 12'd4095;
            12'd3830: PAGE <= 12'd4095;
            12'd3831: PAGE <= 12'd4095;
            12'd3832: PAGE <= 12'd4095;
            12'd3833: PAGE <= 12'd4095;
            12'd3834: PAGE <= 12'd4095;
            12'd3835: PAGE <= 12'd4095;
            12'd3836: PAGE <= 12'd4095;
            12'd3837: PAGE <= 12'd4095;
            12'd3838: PAGE <= 12'd4095;
            12'd3839: PAGE <= 12'd4095;
            12'd3840: PAGE <= 12'd4095;
            12'd3841: PAGE <= 12'd4095;
            12'd3842: PAGE <= 12'd4095;
            12'd3843: PAGE <= 12'd4095;
            12'd3844: PAGE <= 12'd4095;
            12'd3845: PAGE <= 12'd4095;
            12'd3846: PAGE <= 12'd4095;
            12'd3847: PAGE <= 12'd4095;
            12'd3848: PAGE <= 12'd4095;
            12'd3849: PAGE <= 12'd4095;
            12'd3850: PAGE <= 12'd4095;
            12'd3851: PAGE <= 12'd4095;
            12'd3852: PAGE <= 12'd4095;
            12'd3853: PAGE <= 12'd4095;
            12'd3854: PAGE <= 12'd4095;
            12'd3855: PAGE <= 12'd4095;
            12'd3856: PAGE <= 12'd4095;
            12'd3857: PAGE <= 12'd4095;
            12'd3858: PAGE <= 12'd4095;
            12'd3859: PAGE <= 12'd4095;
            12'd3860: PAGE <= 12'd4095;
            12'd3861: PAGE <= 12'd4095;
            12'd3862: PAGE <= 12'd4095;
            12'd3863: PAGE <= 12'd4095;
            12'd3864: PAGE <= 12'd4095;
            12'd3865: PAGE <= 12'd4095;
            12'd3866: PAGE <= 12'd4095;
            12'd3867: PAGE <= 12'd4095;
            12'd3868: PAGE <= 12'd4095;
            12'd3869: PAGE <= 12'd4095;
            12'd3870: PAGE <= 12'd4095;
            12'd3871: PAGE <= 12'd4095;
            12'd3872: PAGE <= 12'd4095;
            12'd3873: PAGE <= 12'd4095;
            12'd3874: PAGE <= 12'd4095;
            12'd3875: PAGE <= 12'd4095;
            12'd3876: PAGE <= 12'd4095;
            12'd3877: PAGE <= 12'd4095;
            12'd3878: PAGE <= 12'd4095;
            12'd3879: PAGE <= 12'd4095;
            12'd3880: PAGE <= 12'd4095;
            12'd3881: PAGE <= 12'd4095;
            12'd3882: PAGE <= 12'd4095;
            12'd3883: PAGE <= 12'd4095;
            12'd3884: PAGE <= 12'd4095;
            12'd3885: PAGE <= 12'd4095;
            12'd3886: PAGE <= 12'd4095;
            12'd3887: PAGE <= 12'd4095;
            12'd3888: PAGE <= 12'd4095;
            12'd3889: PAGE <= 12'd4095;
            12'd3890: PAGE <= 12'd4095;
            12'd3891: PAGE <= 12'd4095;
            12'd3892: PAGE <= 12'd4095;
            12'd3893: PAGE <= 12'd4095;
            12'd3894: PAGE <= 12'd4095;
            12'd3895: PAGE <= 12'd4095;
            12'd3896: PAGE <= 12'd4095;
            12'd3897: PAGE <= 12'd4095;
            12'd3898: PAGE <= 12'd4095;
            12'd3899: PAGE <= 12'd4095;
            12'd3900: PAGE <= 12'd4095;
            12'd3901: PAGE <= 12'd4095;
            12'd3902: PAGE <= 12'd4095;
            12'd3903: PAGE <= 12'd4095;
            12'd3904: PAGE <= 12'd4095;
            12'd3905: PAGE <= 12'd4095;
            12'd3906: PAGE <= 12'd4095;
            12'd3907: PAGE <= 12'd4095;
            12'd3908: PAGE <= 12'd4095;
            12'd3909: PAGE <= 12'd4095;
            12'd3910: PAGE <= 12'd4095;
            12'd3911: PAGE <= 12'd4095;
            12'd3912: PAGE <= 12'd4095;
            12'd3913: PAGE <= 12'd4095;
            12'd3914: PAGE <= 12'd4095;
            12'd3915: PAGE <= 12'd4095;
            12'd3916: PAGE <= 12'd4095;
            12'd3917: PAGE <= 12'd4095;
            12'd3918: PAGE <= 12'd4095;
            12'd3919: PAGE <= 12'd4095;
            12'd3920: PAGE <= 12'd4095;
            12'd3921: PAGE <= 12'd4095;
            12'd3922: PAGE <= 12'd4095;
            12'd3923: PAGE <= 12'd4095;
            12'd3924: PAGE <= 12'd4095;
            12'd3925: PAGE <= 12'd4095;
            12'd3926: PAGE <= 12'd4095;
            12'd3927: PAGE <= 12'd4095;
            12'd3928: PAGE <= 12'd4095;
            12'd3929: PAGE <= 12'd4095;
            12'd3930: PAGE <= 12'd4095;
            12'd3931: PAGE <= 12'd4095;
            12'd3932: PAGE <= 12'd4095;
            12'd3933: PAGE <= 12'd4095;
            12'd3934: PAGE <= 12'd4095;
            12'd3935: PAGE <= 12'd4095;
            12'd3936: PAGE <= 12'd4095;
            12'd3937: PAGE <= 12'd4095;
            12'd3938: PAGE <= 12'd4095;
            12'd3939: PAGE <= 12'd4095;
            12'd3940: PAGE <= 12'd4095;
            12'd3941: PAGE <= 12'd4095;
            12'd3942: PAGE <= 12'd4095;
            12'd3943: PAGE <= 12'd4095;
            12'd3944: PAGE <= 12'd4095;
            12'd3945: PAGE <= 12'd4095;
            12'd3946: PAGE <= 12'd4095;
            12'd3947: PAGE <= 12'd4095;
            12'd3948: PAGE <= 12'd4095;
            12'd3949: PAGE <= 12'd4095;
            12'd3950: PAGE <= 12'd4095;
            12'd3951: PAGE <= 12'd4095;
            12'd3952: PAGE <= 12'd4095;
            12'd3953: PAGE <= 12'd4095;
            12'd3954: PAGE <= 12'd4095;
            12'd3955: PAGE <= 12'd4095;
            12'd3956: PAGE <= 12'd4095;
            12'd3957: PAGE <= 12'd4095;
            12'd3958: PAGE <= 12'd4095;
            12'd3959: PAGE <= 12'd4095;
            12'd3960: PAGE <= 12'd4095;
            12'd3961: PAGE <= 12'd4095;
            12'd3962: PAGE <= 12'd4095;
            12'd3963: PAGE <= 12'd4095;
            12'd3964: PAGE <= 12'd4095;
            12'd3965: PAGE <= 12'd4095;
            12'd3966: PAGE <= 12'd4095;
            12'd3967: PAGE <= 12'd4095;
            12'd3968: PAGE <= 12'd4095;
            12'd3969: PAGE <= 12'd4095;
            12'd3970: PAGE <= 12'd4095;
            12'd3971: PAGE <= 12'd4095;
            12'd3972: PAGE <= 12'd4095;
            12'd3973: PAGE <= 12'd4095;
            12'd3974: PAGE <= 12'd4095;
            12'd3975: PAGE <= 12'd4095;
            12'd3976: PAGE <= 12'd4095;
            12'd3977: PAGE <= 12'd4095;
            12'd3978: PAGE <= 12'd4095;
            12'd3979: PAGE <= 12'd4095;
            12'd3980: PAGE <= 12'd4095;
            12'd3981: PAGE <= 12'd4095;
            12'd3982: PAGE <= 12'd4095;
            12'd3983: PAGE <= 12'd4095;
            12'd3984: PAGE <= 12'd4095;
            12'd3985: PAGE <= 12'd4095;
            12'd3986: PAGE <= 12'd4095;
            12'd3987: PAGE <= 12'd4095;
            12'd3988: PAGE <= 12'd4095;
            12'd3989: PAGE <= 12'd4095;
            12'd3990: PAGE <= 12'd4095;
            12'd3991: PAGE <= 12'd4095;
            12'd3992: PAGE <= 12'd4095;
            12'd3993: PAGE <= 12'd4095;
            12'd3994: PAGE <= 12'd4095;
            12'd3995: PAGE <= 12'd4095;
            12'd3996: PAGE <= 12'd4095;
            12'd3997: PAGE <= 12'd4095;
            12'd3998: PAGE <= 12'd4095;
            12'd3999: PAGE <= 12'd4095;
            12'd4000: PAGE <= 12'd4095;
            12'd4001: PAGE <= 12'd4095;
            12'd4002: PAGE <= 12'd4095;
            12'd4003: PAGE <= 12'd4095;
            12'd4004: PAGE <= 12'd4095;
            12'd4005: PAGE <= 12'd4095;
            12'd4006: PAGE <= 12'd4095;
            12'd4007: PAGE <= 12'd4095;
            12'd4008: PAGE <= 12'd4095;
            12'd4009: PAGE <= 12'd4095;
            12'd4010: PAGE <= 12'd4095;
            12'd4011: PAGE <= 12'd4095;
            12'd4012: PAGE <= 12'd4095;
            12'd4013: PAGE <= 12'd4095;
            12'd4014: PAGE <= 12'd4095;
            12'd4015: PAGE <= 12'd4095;
            12'd4016: PAGE <= 12'd4095;
            12'd4017: PAGE <= 12'd4095;
            12'd4018: PAGE <= 12'd4095;
            12'd4019: PAGE <= 12'd4095;
            12'd4020: PAGE <= 12'd4095;
            12'd4021: PAGE <= 12'd4095;
            12'd4022: PAGE <= 12'd4095;
            12'd4023: PAGE <= 12'd4095;
            12'd4024: PAGE <= 12'd4095;
            12'd4025: PAGE <= 12'd4095;
            12'd4026: PAGE <= 12'd4095;
            12'd4027: PAGE <= 12'd4095;
            12'd4028: PAGE <= 12'd4095;
            12'd4029: PAGE <= 12'd4095;
            12'd4030: PAGE <= 12'd4095;
            12'd4031: PAGE <= 12'd4095;
            12'd4032: PAGE <= 12'd4095;
            12'd4033: PAGE <= 12'd4095;
            12'd4034: PAGE <= 12'd4095;
            12'd4035: PAGE <= 12'd4095;
            12'd4036: PAGE <= 12'd4095;
            12'd4037: PAGE <= 12'd4095;
            12'd4038: PAGE <= 12'd4095;
            12'd4039: PAGE <= 12'd4095;
            12'd4040: PAGE <= 12'd4095;
            12'd4041: PAGE <= 12'd4095;
            12'd4042: PAGE <= 12'd4095;
            12'd4043: PAGE <= 12'd4095;
            12'd4044: PAGE <= 12'd4095;
            12'd4045: PAGE <= 12'd4095;
            12'd4046: PAGE <= 12'd4095;
            12'd4047: PAGE <= 12'd4095;
            12'd4048: PAGE <= 12'd4095;
            12'd4049: PAGE <= 12'd4095;
            12'd4050: PAGE <= 12'd4095;
            12'd4051: PAGE <= 12'd4095;
            12'd4052: PAGE <= 12'd4095;
            12'd4053: PAGE <= 12'd4095;
            12'd4054: PAGE <= 12'd4095;
            12'd4055: PAGE <= 12'd4095;
            12'd4056: PAGE <= 12'd4095;
            12'd4057: PAGE <= 12'd4095;
            12'd4058: PAGE <= 12'd4095;
            12'd4059: PAGE <= 12'd4095;
            12'd4060: PAGE <= 12'd4095;
            12'd4061: PAGE <= 12'd4095;
            12'd4062: PAGE <= 12'd4095;
            12'd4063: PAGE <= 12'd4095;
            12'd4064: PAGE <= 12'd4095;
            12'd4065: PAGE <= 12'd4095;
            12'd4066: PAGE <= 12'd4095;
            12'd4067: PAGE <= 12'd4095;
            12'd4068: PAGE <= 12'd4095;
            12'd4069: PAGE <= 12'd4095;
            12'd4070: PAGE <= 12'd4095;
            12'd4071: PAGE <= 12'd4095;
            12'd4072: PAGE <= 12'd4095;
            12'd4073: PAGE <= 12'd4095;
            12'd4074: PAGE <= 12'd4095;
            12'd4075: PAGE <= 12'd4095;
            12'd4076: PAGE <= 12'd4095;
            12'd4077: PAGE <= 12'd4095;
            12'd4078: PAGE <= 12'd4095;
            12'd4079: PAGE <= 12'd4095;
            12'd4080: PAGE <= 12'd4095;
            12'd4081: PAGE <= 12'd4095;
            12'd4082: PAGE <= 12'd4095;
            12'd4083: PAGE <= 12'd4095;
            12'd4084: PAGE <= 12'd4095;
            12'd4085: PAGE <= 12'd4095;
            12'd4086: PAGE <= 12'd4095;
            12'd4087: PAGE <= 12'd4095;
            12'd4088: PAGE <= 12'd4095;
            12'd4089: PAGE <= 12'd4095;
            12'd4090: PAGE <= 12'd4095;
            12'd4091: PAGE <= 12'd4095;
            12'd4092: PAGE <= 12'd4095;
            12'd4093: PAGE <= 12'd4095;
            12'd4094: PAGE <= 12'd4095;
            12'd4095: PAGE <= 12'd4095;
        endcase
    end
endmodule
