module RelativePageConverter 
(
    input   wire            MCLK,
    input   wire            nCONV,
    input   wire    [11:0]  ABSPAGE,
    output  reg     [11:0]  RELPAGE = 12'd4095
);

always @ (posedge MCLK)
begin
    if(nCONV == 1'b0)
    begin
        case (ABSPAGE)
            12'd0: RELPAGE <= 12'd1862;
            12'd1: RELPAGE <= 12'd331;
            12'd2: RELPAGE <= 12'd853;
            12'd3: RELPAGE <= 12'd1375;
            12'd4: RELPAGE <= 12'd1897;
            12'd5: RELPAGE <= 12'd366;
            12'd6: RELPAGE <= 12'd888;
            12'd7: RELPAGE <= 12'd1410;
            12'd8: RELPAGE <= 12'd1932;
            12'd9: RELPAGE <= 12'd401;
            12'd10: RELPAGE <= 12'd923;
            12'd11: RELPAGE <= 12'd1445;
            12'd12: RELPAGE <= 12'd1967;
            12'd13: RELPAGE <= 12'd436;
            12'd14: RELPAGE <= 12'd958;
            12'd15: RELPAGE <= 12'd1480;
            12'd16: RELPAGE <= 12'd2002;
            12'd17: RELPAGE <= 12'd471;
            12'd18: RELPAGE <= 12'd993;
            12'd19: RELPAGE <= 12'd1515;
            12'd20: RELPAGE <= 12'd2037;
            12'd21: RELPAGE <= 12'd506;
            12'd22: RELPAGE <= 12'd1028;
            12'd23: RELPAGE <= 12'd1550;
            12'd24: RELPAGE <= 12'd19;
            12'd25: RELPAGE <= 12'd541;
            12'd26: RELPAGE <= 12'd1063;
            12'd27: RELPAGE <= 12'd1585;
            12'd28: RELPAGE <= 12'd54;
            12'd29: RELPAGE <= 12'd576;
            12'd30: RELPAGE <= 12'd1098;
            12'd31: RELPAGE <= 12'd1620;
            12'd32: RELPAGE <= 12'd89;
            12'd33: RELPAGE <= 12'd611;
            12'd34: RELPAGE <= 12'd1133;
            12'd35: RELPAGE <= 12'd1655;
            12'd36: RELPAGE <= 12'd124;
            12'd37: RELPAGE <= 12'd646;
            12'd38: RELPAGE <= 12'd1168;
            12'd39: RELPAGE <= 12'd1690;
            12'd40: RELPAGE <= 12'd159;
            12'd41: RELPAGE <= 12'd681;
            12'd42: RELPAGE <= 12'd1203;
            12'd43: RELPAGE <= 12'd1725;
            12'd44: RELPAGE <= 12'd194;
            12'd45: RELPAGE <= 12'd716;
            12'd46: RELPAGE <= 12'd1238;
            12'd47: RELPAGE <= 12'd1760;
            12'd48: RELPAGE <= 12'd229;
            12'd49: RELPAGE <= 12'd751;
            12'd50: RELPAGE <= 12'd1273;
            12'd51: RELPAGE <= 12'd1795;
            12'd52: RELPAGE <= 12'd264;
            12'd53: RELPAGE <= 12'd786;
            12'd54: RELPAGE <= 12'd1308;
            12'd55: RELPAGE <= 12'd1830;
            12'd56: RELPAGE <= 12'd299;
            12'd57: RELPAGE <= 12'd821;
            12'd58: RELPAGE <= 12'd1343;
            12'd59: RELPAGE <= 12'd1865;
            12'd60: RELPAGE <= 12'd334;
            12'd61: RELPAGE <= 12'd856;
            12'd62: RELPAGE <= 12'd1378;
            12'd63: RELPAGE <= 12'd1900;
            12'd64: RELPAGE <= 12'd369;
            12'd65: RELPAGE <= 12'd891;
            12'd66: RELPAGE <= 12'd1413;
            12'd67: RELPAGE <= 12'd1935;
            12'd68: RELPAGE <= 12'd404;
            12'd69: RELPAGE <= 12'd926;
            12'd70: RELPAGE <= 12'd1448;
            12'd71: RELPAGE <= 12'd1970;
            12'd72: RELPAGE <= 12'd439;
            12'd73: RELPAGE <= 12'd961;
            12'd74: RELPAGE <= 12'd1483;
            12'd75: RELPAGE <= 12'd2005;
            12'd76: RELPAGE <= 12'd474;
            12'd77: RELPAGE <= 12'd996;
            12'd78: RELPAGE <= 12'd1518;
            12'd79: RELPAGE <= 12'd2040;
            12'd80: RELPAGE <= 12'd509;
            12'd81: RELPAGE <= 12'd1031;
            12'd82: RELPAGE <= 12'd1553;
            12'd83: RELPAGE <= 12'd22;
            12'd84: RELPAGE <= 12'd544;
            12'd85: RELPAGE <= 12'd1066;
            12'd86: RELPAGE <= 12'd1588;
            12'd87: RELPAGE <= 12'd57;
            12'd88: RELPAGE <= 12'd579;
            12'd89: RELPAGE <= 12'd1101;
            12'd90: RELPAGE <= 12'd1623;
            12'd91: RELPAGE <= 12'd92;
            12'd92: RELPAGE <= 12'd614;
            12'd93: RELPAGE <= 12'd1136;
            12'd94: RELPAGE <= 12'd1658;
            12'd95: RELPAGE <= 12'd127;
            12'd96: RELPAGE <= 12'd649;
            12'd97: RELPAGE <= 12'd1171;
            12'd98: RELPAGE <= 12'd1693;
            12'd99: RELPAGE <= 12'd162;
            12'd100: RELPAGE <= 12'd684;
            12'd101: RELPAGE <= 12'd1206;
            12'd102: RELPAGE <= 12'd1728;
            12'd103: RELPAGE <= 12'd197;
            12'd104: RELPAGE <= 12'd719;
            12'd105: RELPAGE <= 12'd1241;
            12'd106: RELPAGE <= 12'd1763;
            12'd107: RELPAGE <= 12'd232;
            12'd108: RELPAGE <= 12'd754;
            12'd109: RELPAGE <= 12'd1276;
            12'd110: RELPAGE <= 12'd1798;
            12'd111: RELPAGE <= 12'd267;
            12'd112: RELPAGE <= 12'd789;
            12'd113: RELPAGE <= 12'd1311;
            12'd114: RELPAGE <= 12'd1833;
            12'd115: RELPAGE <= 12'd302;
            12'd116: RELPAGE <= 12'd824;
            12'd117: RELPAGE <= 12'd1346;
            12'd118: RELPAGE <= 12'd1868;
            12'd119: RELPAGE <= 12'd337;
            12'd120: RELPAGE <= 12'd859;
            12'd121: RELPAGE <= 12'd1381;
            12'd122: RELPAGE <= 12'd1903;
            12'd123: RELPAGE <= 12'd372;
            12'd124: RELPAGE <= 12'd894;
            12'd125: RELPAGE <= 12'd1416;
            12'd126: RELPAGE <= 12'd1938;
            12'd127: RELPAGE <= 12'd407;
            12'd128: RELPAGE <= 12'd929;
            12'd129: RELPAGE <= 12'd1451;
            12'd130: RELPAGE <= 12'd1973;
            12'd131: RELPAGE <= 12'd442;
            12'd132: RELPAGE <= 12'd964;
            12'd133: RELPAGE <= 12'd1486;
            12'd134: RELPAGE <= 12'd2008;
            12'd135: RELPAGE <= 12'd477;
            12'd136: RELPAGE <= 12'd999;
            12'd137: RELPAGE <= 12'd1521;
            12'd138: RELPAGE <= 12'd2043;
            12'd139: RELPAGE <= 12'd512;
            12'd140: RELPAGE <= 12'd1034;
            12'd141: RELPAGE <= 12'd1556;
            12'd142: RELPAGE <= 12'd25;
            12'd143: RELPAGE <= 12'd547;
            12'd144: RELPAGE <= 12'd1069;
            12'd145: RELPAGE <= 12'd1591;
            12'd146: RELPAGE <= 12'd60;
            12'd147: RELPAGE <= 12'd582;
            12'd148: RELPAGE <= 12'd1104;
            12'd149: RELPAGE <= 12'd1626;
            12'd150: RELPAGE <= 12'd95;
            12'd151: RELPAGE <= 12'd617;
            12'd152: RELPAGE <= 12'd1139;
            12'd153: RELPAGE <= 12'd1661;
            12'd154: RELPAGE <= 12'd130;
            12'd155: RELPAGE <= 12'd652;
            12'd156: RELPAGE <= 12'd1174;
            12'd157: RELPAGE <= 12'd1696;
            12'd158: RELPAGE <= 12'd165;
            12'd159: RELPAGE <= 12'd687;
            12'd160: RELPAGE <= 12'd1209;
            12'd161: RELPAGE <= 12'd1731;
            12'd162: RELPAGE <= 12'd200;
            12'd163: RELPAGE <= 12'd722;
            12'd164: RELPAGE <= 12'd1244;
            12'd165: RELPAGE <= 12'd1766;
            12'd166: RELPAGE <= 12'd235;
            12'd167: RELPAGE <= 12'd757;
            12'd168: RELPAGE <= 12'd1279;
            12'd169: RELPAGE <= 12'd1801;
            12'd170: RELPAGE <= 12'd270;
            12'd171: RELPAGE <= 12'd792;
            12'd172: RELPAGE <= 12'd1314;
            12'd173: RELPAGE <= 12'd1836;
            12'd174: RELPAGE <= 12'd305;
            12'd175: RELPAGE <= 12'd827;
            12'd176: RELPAGE <= 12'd1349;
            12'd177: RELPAGE <= 12'd1871;
            12'd178: RELPAGE <= 12'd340;
            12'd179: RELPAGE <= 12'd862;
            12'd180: RELPAGE <= 12'd1384;
            12'd181: RELPAGE <= 12'd1906;
            12'd182: RELPAGE <= 12'd375;
            12'd183: RELPAGE <= 12'd897;
            12'd184: RELPAGE <= 12'd1419;
            12'd185: RELPAGE <= 12'd1941;
            12'd186: RELPAGE <= 12'd410;
            12'd187: RELPAGE <= 12'd932;
            12'd188: RELPAGE <= 12'd1454;
            12'd189: RELPAGE <= 12'd1976;
            12'd190: RELPAGE <= 12'd445;
            12'd191: RELPAGE <= 12'd967;
            12'd192: RELPAGE <= 12'd1489;
            12'd193: RELPAGE <= 12'd2011;
            12'd194: RELPAGE <= 12'd480;
            12'd195: RELPAGE <= 12'd1002;
            12'd196: RELPAGE <= 12'd1524;
            12'd197: RELPAGE <= 12'd2046;
            12'd198: RELPAGE <= 12'd515;
            12'd199: RELPAGE <= 12'd1037;
            12'd200: RELPAGE <= 12'd1559;
            12'd201: RELPAGE <= 12'd28;
            12'd202: RELPAGE <= 12'd550;
            12'd203: RELPAGE <= 12'd1072;
            12'd204: RELPAGE <= 12'd1594;
            12'd205: RELPAGE <= 12'd63;
            12'd206: RELPAGE <= 12'd585;
            12'd207: RELPAGE <= 12'd1107;
            12'd208: RELPAGE <= 12'd1629;
            12'd209: RELPAGE <= 12'd98;
            12'd210: RELPAGE <= 12'd620;
            12'd211: RELPAGE <= 12'd1142;
            12'd212: RELPAGE <= 12'd1664;
            12'd213: RELPAGE <= 12'd133;
            12'd214: RELPAGE <= 12'd655;
            12'd215: RELPAGE <= 12'd1177;
            12'd216: RELPAGE <= 12'd1699;
            12'd217: RELPAGE <= 12'd168;
            12'd218: RELPAGE <= 12'd690;
            12'd219: RELPAGE <= 12'd1212;
            12'd220: RELPAGE <= 12'd1734;
            12'd221: RELPAGE <= 12'd203;
            12'd222: RELPAGE <= 12'd725;
            12'd223: RELPAGE <= 12'd1247;
            12'd224: RELPAGE <= 12'd1769;
            12'd225: RELPAGE <= 12'd238;
            12'd226: RELPAGE <= 12'd760;
            12'd227: RELPAGE <= 12'd1282;
            12'd228: RELPAGE <= 12'd1804;
            12'd229: RELPAGE <= 12'd273;
            12'd230: RELPAGE <= 12'd795;
            12'd231: RELPAGE <= 12'd1317;
            12'd232: RELPAGE <= 12'd1839;
            12'd233: RELPAGE <= 12'd308;
            12'd234: RELPAGE <= 12'd830;
            12'd235: RELPAGE <= 12'd1352;
            12'd236: RELPAGE <= 12'd1874;
            12'd237: RELPAGE <= 12'd343;
            12'd238: RELPAGE <= 12'd865;
            12'd239: RELPAGE <= 12'd1387;
            12'd240: RELPAGE <= 12'd1909;
            12'd241: RELPAGE <= 12'd378;
            12'd242: RELPAGE <= 12'd900;
            12'd243: RELPAGE <= 12'd1422;
            12'd244: RELPAGE <= 12'd1944;
            12'd245: RELPAGE <= 12'd413;
            12'd246: RELPAGE <= 12'd935;
            12'd247: RELPAGE <= 12'd1457;
            12'd248: RELPAGE <= 12'd1979;
            12'd249: RELPAGE <= 12'd448;
            12'd250: RELPAGE <= 12'd970;
            12'd251: RELPAGE <= 12'd1492;
            12'd252: RELPAGE <= 12'd2014;
            12'd253: RELPAGE <= 12'd483;
            12'd254: RELPAGE <= 12'd1005;
            12'd255: RELPAGE <= 12'd1527;
            12'd256: RELPAGE <= 12'd2049;
            12'd257: RELPAGE <= 12'd518;
            12'd258: RELPAGE <= 12'd1040;
            12'd259: RELPAGE <= 12'd1562;
            12'd260: RELPAGE <= 12'd31;
            12'd261: RELPAGE <= 12'd553;
            12'd262: RELPAGE <= 12'd1075;
            12'd263: RELPAGE <= 12'd1597;
            12'd264: RELPAGE <= 12'd66;
            12'd265: RELPAGE <= 12'd588;
            12'd266: RELPAGE <= 12'd1110;
            12'd267: RELPAGE <= 12'd1632;
            12'd268: RELPAGE <= 12'd101;
            12'd269: RELPAGE <= 12'd623;
            12'd270: RELPAGE <= 12'd1145;
            12'd271: RELPAGE <= 12'd1667;
            12'd272: RELPAGE <= 12'd136;
            12'd273: RELPAGE <= 12'd658;
            12'd274: RELPAGE <= 12'd1180;
            12'd275: RELPAGE <= 12'd1702;
            12'd276: RELPAGE <= 12'd171;
            12'd277: RELPAGE <= 12'd693;
            12'd278: RELPAGE <= 12'd1215;
            12'd279: RELPAGE <= 12'd1737;
            12'd280: RELPAGE <= 12'd206;
            12'd281: RELPAGE <= 12'd728;
            12'd282: RELPAGE <= 12'd1250;
            12'd283: RELPAGE <= 12'd1772;
            12'd284: RELPAGE <= 12'd241;
            12'd285: RELPAGE <= 12'd763;
            12'd286: RELPAGE <= 12'd1285;
            12'd287: RELPAGE <= 12'd1807;
            12'd288: RELPAGE <= 12'd276;
            12'd289: RELPAGE <= 12'd798;
            12'd290: RELPAGE <= 12'd1320;
            12'd291: RELPAGE <= 12'd1842;
            12'd292: RELPAGE <= 12'd311;
            12'd293: RELPAGE <= 12'd833;
            12'd294: RELPAGE <= 12'd1355;
            12'd295: RELPAGE <= 12'd1877;
            12'd296: RELPAGE <= 12'd346;
            12'd297: RELPAGE <= 12'd868;
            12'd298: RELPAGE <= 12'd1390;
            12'd299: RELPAGE <= 12'd1912;
            12'd300: RELPAGE <= 12'd381;
            12'd301: RELPAGE <= 12'd903;
            12'd302: RELPAGE <= 12'd1425;
            12'd303: RELPAGE <= 12'd1947;
            12'd304: RELPAGE <= 12'd416;
            12'd305: RELPAGE <= 12'd938;
            12'd306: RELPAGE <= 12'd1460;
            12'd307: RELPAGE <= 12'd1982;
            12'd308: RELPAGE <= 12'd451;
            12'd309: RELPAGE <= 12'd973;
            12'd310: RELPAGE <= 12'd1495;
            12'd311: RELPAGE <= 12'd2017;
            12'd312: RELPAGE <= 12'd486;
            12'd313: RELPAGE <= 12'd1008;
            12'd314: RELPAGE <= 12'd1530;
            12'd315: RELPAGE <= 12'd2052;
            12'd316: RELPAGE <= 12'd521;
            12'd317: RELPAGE <= 12'd1043;
            12'd318: RELPAGE <= 12'd1565;
            12'd319: RELPAGE <= 12'd34;
            12'd320: RELPAGE <= 12'd556;
            12'd321: RELPAGE <= 12'd1078;
            12'd322: RELPAGE <= 12'd1600;
            12'd323: RELPAGE <= 12'd69;
            12'd324: RELPAGE <= 12'd591;
            12'd325: RELPAGE <= 12'd1113;
            12'd326: RELPAGE <= 12'd1635;
            12'd327: RELPAGE <= 12'd104;
            12'd328: RELPAGE <= 12'd626;
            12'd329: RELPAGE <= 12'd1148;
            12'd330: RELPAGE <= 12'd1670;
            12'd331: RELPAGE <= 12'd139;
            12'd332: RELPAGE <= 12'd661;
            12'd333: RELPAGE <= 12'd1183;
            12'd334: RELPAGE <= 12'd1705;
            12'd335: RELPAGE <= 12'd174;
            12'd336: RELPAGE <= 12'd696;
            12'd337: RELPAGE <= 12'd1218;
            12'd338: RELPAGE <= 12'd1740;
            12'd339: RELPAGE <= 12'd209;
            12'd340: RELPAGE <= 12'd731;
            12'd341: RELPAGE <= 12'd1253;
            12'd342: RELPAGE <= 12'd1775;
            12'd343: RELPAGE <= 12'd244;
            12'd344: RELPAGE <= 12'd766;
            12'd345: RELPAGE <= 12'd1288;
            12'd346: RELPAGE <= 12'd1810;
            12'd347: RELPAGE <= 12'd279;
            12'd348: RELPAGE <= 12'd801;
            12'd349: RELPAGE <= 12'd1323;
            12'd350: RELPAGE <= 12'd1845;
            12'd351: RELPAGE <= 12'd314;
            12'd352: RELPAGE <= 12'd836;
            12'd353: RELPAGE <= 12'd1358;
            12'd354: RELPAGE <= 12'd1880;
            12'd355: RELPAGE <= 12'd349;
            12'd356: RELPAGE <= 12'd871;
            12'd357: RELPAGE <= 12'd1393;
            12'd358: RELPAGE <= 12'd1915;
            12'd359: RELPAGE <= 12'd384;
            12'd360: RELPAGE <= 12'd906;
            12'd361: RELPAGE <= 12'd1428;
            12'd362: RELPAGE <= 12'd1950;
            12'd363: RELPAGE <= 12'd419;
            12'd364: RELPAGE <= 12'd941;
            12'd365: RELPAGE <= 12'd1463;
            12'd366: RELPAGE <= 12'd1985;
            12'd367: RELPAGE <= 12'd454;
            12'd368: RELPAGE <= 12'd976;
            12'd369: RELPAGE <= 12'd1498;
            12'd370: RELPAGE <= 12'd2020;
            12'd371: RELPAGE <= 12'd489;
            12'd372: RELPAGE <= 12'd1011;
            12'd373: RELPAGE <= 12'd1533;
            12'd374: RELPAGE <= 12'd2;
            12'd375: RELPAGE <= 12'd524;
            12'd376: RELPAGE <= 12'd1046;
            12'd377: RELPAGE <= 12'd1568;
            12'd378: RELPAGE <= 12'd37;
            12'd379: RELPAGE <= 12'd559;
            12'd380: RELPAGE <= 12'd1081;
            12'd381: RELPAGE <= 12'd1603;
            12'd382: RELPAGE <= 12'd72;
            12'd383: RELPAGE <= 12'd594;
            12'd384: RELPAGE <= 12'd1116;
            12'd385: RELPAGE <= 12'd1638;
            12'd386: RELPAGE <= 12'd107;
            12'd387: RELPAGE <= 12'd629;
            12'd388: RELPAGE <= 12'd1151;
            12'd389: RELPAGE <= 12'd1673;
            12'd390: RELPAGE <= 12'd142;
            12'd391: RELPAGE <= 12'd664;
            12'd392: RELPAGE <= 12'd1186;
            12'd393: RELPAGE <= 12'd1708;
            12'd394: RELPAGE <= 12'd177;
            12'd395: RELPAGE <= 12'd699;
            12'd396: RELPAGE <= 12'd1221;
            12'd397: RELPAGE <= 12'd1743;
            12'd398: RELPAGE <= 12'd212;
            12'd399: RELPAGE <= 12'd734;
            12'd400: RELPAGE <= 12'd1256;
            12'd401: RELPAGE <= 12'd1778;
            12'd402: RELPAGE <= 12'd247;
            12'd403: RELPAGE <= 12'd769;
            12'd404: RELPAGE <= 12'd1291;
            12'd405: RELPAGE <= 12'd1813;
            12'd406: RELPAGE <= 12'd282;
            12'd407: RELPAGE <= 12'd804;
            12'd408: RELPAGE <= 12'd1326;
            12'd409: RELPAGE <= 12'd1848;
            12'd410: RELPAGE <= 12'd317;
            12'd411: RELPAGE <= 12'd839;
            12'd412: RELPAGE <= 12'd1361;
            12'd413: RELPAGE <= 12'd1883;
            12'd414: RELPAGE <= 12'd352;
            12'd415: RELPAGE <= 12'd874;
            12'd416: RELPAGE <= 12'd1396;
            12'd417: RELPAGE <= 12'd1918;
            12'd418: RELPAGE <= 12'd387;
            12'd419: RELPAGE <= 12'd909;
            12'd420: RELPAGE <= 12'd1431;
            12'd421: RELPAGE <= 12'd1953;
            12'd422: RELPAGE <= 12'd422;
            12'd423: RELPAGE <= 12'd944;
            12'd424: RELPAGE <= 12'd1466;
            12'd425: RELPAGE <= 12'd1988;
            12'd426: RELPAGE <= 12'd457;
            12'd427: RELPAGE <= 12'd979;
            12'd428: RELPAGE <= 12'd1501;
            12'd429: RELPAGE <= 12'd2023;
            12'd430: RELPAGE <= 12'd492;
            12'd431: RELPAGE <= 12'd1014;
            12'd432: RELPAGE <= 12'd1536;
            12'd433: RELPAGE <= 12'd5;
            12'd434: RELPAGE <= 12'd527;
            12'd435: RELPAGE <= 12'd1049;
            12'd436: RELPAGE <= 12'd1571;
            12'd437: RELPAGE <= 12'd40;
            12'd438: RELPAGE <= 12'd562;
            12'd439: RELPAGE <= 12'd1084;
            12'd440: RELPAGE <= 12'd1606;
            12'd441: RELPAGE <= 12'd75;
            12'd442: RELPAGE <= 12'd597;
            12'd443: RELPAGE <= 12'd1119;
            12'd444: RELPAGE <= 12'd1641;
            12'd445: RELPAGE <= 12'd110;
            12'd446: RELPAGE <= 12'd632;
            12'd447: RELPAGE <= 12'd1154;
            12'd448: RELPAGE <= 12'd1676;
            12'd449: RELPAGE <= 12'd145;
            12'd450: RELPAGE <= 12'd667;
            12'd451: RELPAGE <= 12'd1189;
            12'd452: RELPAGE <= 12'd1711;
            12'd453: RELPAGE <= 12'd180;
            12'd454: RELPAGE <= 12'd702;
            12'd455: RELPAGE <= 12'd1224;
            12'd456: RELPAGE <= 12'd1746;
            12'd457: RELPAGE <= 12'd215;
            12'd458: RELPAGE <= 12'd737;
            12'd459: RELPAGE <= 12'd1259;
            12'd460: RELPAGE <= 12'd1781;
            12'd461: RELPAGE <= 12'd250;
            12'd462: RELPAGE <= 12'd772;
            12'd463: RELPAGE <= 12'd1294;
            12'd464: RELPAGE <= 12'd1816;
            12'd465: RELPAGE <= 12'd285;
            12'd466: RELPAGE <= 12'd807;
            12'd467: RELPAGE <= 12'd1329;
            12'd468: RELPAGE <= 12'd1851;
            12'd469: RELPAGE <= 12'd320;
            12'd470: RELPAGE <= 12'd842;
            12'd471: RELPAGE <= 12'd1364;
            12'd472: RELPAGE <= 12'd1886;
            12'd473: RELPAGE <= 12'd355;
            12'd474: RELPAGE <= 12'd877;
            12'd475: RELPAGE <= 12'd1399;
            12'd476: RELPAGE <= 12'd1921;
            12'd477: RELPAGE <= 12'd390;
            12'd478: RELPAGE <= 12'd912;
            12'd479: RELPAGE <= 12'd1434;
            12'd480: RELPAGE <= 12'd1956;
            12'd481: RELPAGE <= 12'd425;
            12'd482: RELPAGE <= 12'd947;
            12'd483: RELPAGE <= 12'd1469;
            12'd484: RELPAGE <= 12'd1991;
            12'd485: RELPAGE <= 12'd460;
            12'd486: RELPAGE <= 12'd982;
            12'd487: RELPAGE <= 12'd1504;
            12'd488: RELPAGE <= 12'd2026;
            12'd489: RELPAGE <= 12'd495;
            12'd490: RELPAGE <= 12'd1017;
            12'd491: RELPAGE <= 12'd1539;
            12'd492: RELPAGE <= 12'd8;
            12'd493: RELPAGE <= 12'd530;
            12'd494: RELPAGE <= 12'd1052;
            12'd495: RELPAGE <= 12'd1574;
            12'd496: RELPAGE <= 12'd43;
            12'd497: RELPAGE <= 12'd565;
            12'd498: RELPAGE <= 12'd1087;
            12'd499: RELPAGE <= 12'd1609;
            12'd500: RELPAGE <= 12'd78;
            12'd501: RELPAGE <= 12'd600;
            12'd502: RELPAGE <= 12'd1122;
            12'd503: RELPAGE <= 12'd1644;
            12'd504: RELPAGE <= 12'd113;
            12'd505: RELPAGE <= 12'd635;
            12'd506: RELPAGE <= 12'd1157;
            12'd507: RELPAGE <= 12'd1679;
            12'd508: RELPAGE <= 12'd148;
            12'd509: RELPAGE <= 12'd670;
            12'd510: RELPAGE <= 12'd1192;
            12'd511: RELPAGE <= 12'd1714;
            12'd512: RELPAGE <= 12'd183;
            12'd513: RELPAGE <= 12'd705;
            12'd514: RELPAGE <= 12'd1227;
            12'd515: RELPAGE <= 12'd1749;
            12'd516: RELPAGE <= 12'd218;
            12'd517: RELPAGE <= 12'd740;
            12'd518: RELPAGE <= 12'd1262;
            12'd519: RELPAGE <= 12'd1784;
            12'd520: RELPAGE <= 12'd253;
            12'd521: RELPAGE <= 12'd775;
            12'd522: RELPAGE <= 12'd1297;
            12'd523: RELPAGE <= 12'd1819;
            12'd524: RELPAGE <= 12'd288;
            12'd525: RELPAGE <= 12'd810;
            12'd526: RELPAGE <= 12'd1332;
            12'd527: RELPAGE <= 12'd1854;
            12'd528: RELPAGE <= 12'd323;
            12'd529: RELPAGE <= 12'd845;
            12'd530: RELPAGE <= 12'd1367;
            12'd531: RELPAGE <= 12'd1889;
            12'd532: RELPAGE <= 12'd358;
            12'd533: RELPAGE <= 12'd880;
            12'd534: RELPAGE <= 12'd1402;
            12'd535: RELPAGE <= 12'd1924;
            12'd536: RELPAGE <= 12'd393;
            12'd537: RELPAGE <= 12'd915;
            12'd538: RELPAGE <= 12'd1437;
            12'd539: RELPAGE <= 12'd1959;
            12'd540: RELPAGE <= 12'd428;
            12'd541: RELPAGE <= 12'd950;
            12'd542: RELPAGE <= 12'd1472;
            12'd543: RELPAGE <= 12'd1994;
            12'd544: RELPAGE <= 12'd463;
            12'd545: RELPAGE <= 12'd985;
            12'd546: RELPAGE <= 12'd1507;
            12'd547: RELPAGE <= 12'd2029;
            12'd548: RELPAGE <= 12'd498;
            12'd549: RELPAGE <= 12'd1020;
            12'd550: RELPAGE <= 12'd1542;
            12'd551: RELPAGE <= 12'd11;
            12'd552: RELPAGE <= 12'd533;
            12'd553: RELPAGE <= 12'd1055;
            12'd554: RELPAGE <= 12'd1577;
            12'd555: RELPAGE <= 12'd46;
            12'd556: RELPAGE <= 12'd568;
            12'd557: RELPAGE <= 12'd1090;
            12'd558: RELPAGE <= 12'd1612;
            12'd559: RELPAGE <= 12'd81;
            12'd560: RELPAGE <= 12'd603;
            12'd561: RELPAGE <= 12'd1125;
            12'd562: RELPAGE <= 12'd1647;
            12'd563: RELPAGE <= 12'd116;
            12'd564: RELPAGE <= 12'd638;
            12'd565: RELPAGE <= 12'd1160;
            12'd566: RELPAGE <= 12'd1682;
            12'd567: RELPAGE <= 12'd151;
            12'd568: RELPAGE <= 12'd673;
            12'd569: RELPAGE <= 12'd1195;
            12'd570: RELPAGE <= 12'd1717;
            12'd571: RELPAGE <= 12'd186;
            12'd572: RELPAGE <= 12'd708;
            12'd573: RELPAGE <= 12'd1230;
            12'd574: RELPAGE <= 12'd1752;
            12'd575: RELPAGE <= 12'd221;
            12'd576: RELPAGE <= 12'd743;
            12'd577: RELPAGE <= 12'd1265;
            12'd578: RELPAGE <= 12'd1787;
            12'd579: RELPAGE <= 12'd256;
            12'd580: RELPAGE <= 12'd778;
            12'd581: RELPAGE <= 12'd1300;
            12'd582: RELPAGE <= 12'd1822;
            12'd583: RELPAGE <= 12'd291;
            12'd584: RELPAGE <= 12'd813;
            12'd585: RELPAGE <= 12'd1335;
            12'd586: RELPAGE <= 12'd1857;
            12'd587: RELPAGE <= 12'd326;
            12'd588: RELPAGE <= 12'd848;
            12'd589: RELPAGE <= 12'd1370;
            12'd590: RELPAGE <= 12'd1892;
            12'd591: RELPAGE <= 12'd361;
            12'd592: RELPAGE <= 12'd883;
            12'd593: RELPAGE <= 12'd1405;
            12'd594: RELPAGE <= 12'd1927;
            12'd595: RELPAGE <= 12'd396;
            12'd596: RELPAGE <= 12'd918;
            12'd597: RELPAGE <= 12'd1440;
            12'd598: RELPAGE <= 12'd1962;
            12'd599: RELPAGE <= 12'd431;
            12'd600: RELPAGE <= 12'd953;
            12'd601: RELPAGE <= 12'd1475;
            12'd602: RELPAGE <= 12'd1997;
            12'd603: RELPAGE <= 12'd466;
            12'd604: RELPAGE <= 12'd988;
            12'd605: RELPAGE <= 12'd1510;
            12'd606: RELPAGE <= 12'd2032;
            12'd607: RELPAGE <= 12'd501;
            12'd608: RELPAGE <= 12'd1023;
            12'd609: RELPAGE <= 12'd1545;
            12'd610: RELPAGE <= 12'd14;
            12'd611: RELPAGE <= 12'd536;
            12'd612: RELPAGE <= 12'd1058;
            12'd613: RELPAGE <= 12'd1580;
            12'd614: RELPAGE <= 12'd49;
            12'd615: RELPAGE <= 12'd571;
            12'd616: RELPAGE <= 12'd1093;
            12'd617: RELPAGE <= 12'd1615;
            12'd618: RELPAGE <= 12'd84;
            12'd619: RELPAGE <= 12'd606;
            12'd620: RELPAGE <= 12'd1128;
            12'd621: RELPAGE <= 12'd1650;
            12'd622: RELPAGE <= 12'd119;
            12'd623: RELPAGE <= 12'd641;
            12'd624: RELPAGE <= 12'd1163;
            12'd625: RELPAGE <= 12'd1685;
            12'd626: RELPAGE <= 12'd154;
            12'd627: RELPAGE <= 12'd676;
            12'd628: RELPAGE <= 12'd1198;
            12'd629: RELPAGE <= 12'd1720;
            12'd630: RELPAGE <= 12'd189;
            12'd631: RELPAGE <= 12'd711;
            12'd632: RELPAGE <= 12'd1233;
            12'd633: RELPAGE <= 12'd1755;
            12'd634: RELPAGE <= 12'd224;
            12'd635: RELPAGE <= 12'd746;
            12'd636: RELPAGE <= 12'd1268;
            12'd637: RELPAGE <= 12'd1790;
            12'd638: RELPAGE <= 12'd259;
            12'd639: RELPAGE <= 12'd781;
            12'd640: RELPAGE <= 12'd1303;
            12'd641: RELPAGE <= 12'd1825;
            12'd642: RELPAGE <= 12'd294;
            12'd643: RELPAGE <= 12'd816;
            12'd644: RELPAGE <= 12'd1338;
            12'd645: RELPAGE <= 12'd1860;
            12'd646: RELPAGE <= 12'd329;
            12'd647: RELPAGE <= 12'd851;
            12'd648: RELPAGE <= 12'd1373;
            12'd649: RELPAGE <= 12'd1895;
            12'd650: RELPAGE <= 12'd364;
            12'd651: RELPAGE <= 12'd886;
            12'd652: RELPAGE <= 12'd1408;
            12'd653: RELPAGE <= 12'd1930;
            12'd654: RELPAGE <= 12'd399;
            12'd655: RELPAGE <= 12'd921;
            12'd656: RELPAGE <= 12'd1443;
            12'd657: RELPAGE <= 12'd1965;
            12'd658: RELPAGE <= 12'd434;
            12'd659: RELPAGE <= 12'd956;
            12'd660: RELPAGE <= 12'd1478;
            12'd661: RELPAGE <= 12'd2000;
            12'd662: RELPAGE <= 12'd469;
            12'd663: RELPAGE <= 12'd991;
            12'd664: RELPAGE <= 12'd1513;
            12'd665: RELPAGE <= 12'd2035;
            12'd666: RELPAGE <= 12'd504;
            12'd667: RELPAGE <= 12'd1026;
            12'd668: RELPAGE <= 12'd1548;
            12'd669: RELPAGE <= 12'd17;
            12'd670: RELPAGE <= 12'd539;
            12'd671: RELPAGE <= 12'd1061;
            12'd672: RELPAGE <= 12'd1583;
            12'd673: RELPAGE <= 12'd52;
            12'd674: RELPAGE <= 12'd574;
            12'd675: RELPAGE <= 12'd1096;
            12'd676: RELPAGE <= 12'd1618;
            12'd677: RELPAGE <= 12'd87;
            12'd678: RELPAGE <= 12'd609;
            12'd679: RELPAGE <= 12'd1131;
            12'd680: RELPAGE <= 12'd1653;
            12'd681: RELPAGE <= 12'd122;
            12'd682: RELPAGE <= 12'd644;
            12'd683: RELPAGE <= 12'd1166;
            12'd684: RELPAGE <= 12'd1688;
            12'd685: RELPAGE <= 12'd157;
            12'd686: RELPAGE <= 12'd679;
            12'd687: RELPAGE <= 12'd1201;
            12'd688: RELPAGE <= 12'd1723;
            12'd689: RELPAGE <= 12'd192;
            12'd690: RELPAGE <= 12'd714;
            12'd691: RELPAGE <= 12'd1236;
            12'd692: RELPAGE <= 12'd1758;
            12'd693: RELPAGE <= 12'd227;
            12'd694: RELPAGE <= 12'd749;
            12'd695: RELPAGE <= 12'd1271;
            12'd696: RELPAGE <= 12'd1793;
            12'd697: RELPAGE <= 12'd262;
            12'd698: RELPAGE <= 12'd784;
            12'd699: RELPAGE <= 12'd1306;
            12'd700: RELPAGE <= 12'd1828;
            12'd701: RELPAGE <= 12'd297;
            12'd702: RELPAGE <= 12'd819;
            12'd703: RELPAGE <= 12'd1341;
            12'd704: RELPAGE <= 12'd1863;
            12'd705: RELPAGE <= 12'd332;
            12'd706: RELPAGE <= 12'd854;
            12'd707: RELPAGE <= 12'd1376;
            12'd708: RELPAGE <= 12'd1898;
            12'd709: RELPAGE <= 12'd367;
            12'd710: RELPAGE <= 12'd889;
            12'd711: RELPAGE <= 12'd1411;
            12'd712: RELPAGE <= 12'd1933;
            12'd713: RELPAGE <= 12'd402;
            12'd714: RELPAGE <= 12'd924;
            12'd715: RELPAGE <= 12'd1446;
            12'd716: RELPAGE <= 12'd1968;
            12'd717: RELPAGE <= 12'd437;
            12'd718: RELPAGE <= 12'd959;
            12'd719: RELPAGE <= 12'd1481;
            12'd720: RELPAGE <= 12'd2003;
            12'd721: RELPAGE <= 12'd472;
            12'd722: RELPAGE <= 12'd994;
            12'd723: RELPAGE <= 12'd1516;
            12'd724: RELPAGE <= 12'd2038;
            12'd725: RELPAGE <= 12'd507;
            12'd726: RELPAGE <= 12'd1029;
            12'd727: RELPAGE <= 12'd1551;
            12'd728: RELPAGE <= 12'd20;
            12'd729: RELPAGE <= 12'd542;
            12'd730: RELPAGE <= 12'd1064;
            12'd731: RELPAGE <= 12'd1586;
            12'd732: RELPAGE <= 12'd55;
            12'd733: RELPAGE <= 12'd577;
            12'd734: RELPAGE <= 12'd1099;
            12'd735: RELPAGE <= 12'd1621;
            12'd736: RELPAGE <= 12'd90;
            12'd737: RELPAGE <= 12'd612;
            12'd738: RELPAGE <= 12'd1134;
            12'd739: RELPAGE <= 12'd1656;
            12'd740: RELPAGE <= 12'd125;
            12'd741: RELPAGE <= 12'd647;
            12'd742: RELPAGE <= 12'd1169;
            12'd743: RELPAGE <= 12'd1691;
            12'd744: RELPAGE <= 12'd160;
            12'd745: RELPAGE <= 12'd682;
            12'd746: RELPAGE <= 12'd1204;
            12'd747: RELPAGE <= 12'd1726;
            12'd748: RELPAGE <= 12'd195;
            12'd749: RELPAGE <= 12'd717;
            12'd750: RELPAGE <= 12'd1239;
            12'd751: RELPAGE <= 12'd1761;
            12'd752: RELPAGE <= 12'd230;
            12'd753: RELPAGE <= 12'd752;
            12'd754: RELPAGE <= 12'd1274;
            12'd755: RELPAGE <= 12'd1796;
            12'd756: RELPAGE <= 12'd265;
            12'd757: RELPAGE <= 12'd787;
            12'd758: RELPAGE <= 12'd1309;
            12'd759: RELPAGE <= 12'd1831;
            12'd760: RELPAGE <= 12'd300;
            12'd761: RELPAGE <= 12'd822;
            12'd762: RELPAGE <= 12'd1344;
            12'd763: RELPAGE <= 12'd1866;
            12'd764: RELPAGE <= 12'd335;
            12'd765: RELPAGE <= 12'd857;
            12'd766: RELPAGE <= 12'd1379;
            12'd767: RELPAGE <= 12'd1901;
            12'd768: RELPAGE <= 12'd370;
            12'd769: RELPAGE <= 12'd892;
            12'd770: RELPAGE <= 12'd1414;
            12'd771: RELPAGE <= 12'd1936;
            12'd772: RELPAGE <= 12'd405;
            12'd773: RELPAGE <= 12'd927;
            12'd774: RELPAGE <= 12'd1449;
            12'd775: RELPAGE <= 12'd1971;
            12'd776: RELPAGE <= 12'd440;
            12'd777: RELPAGE <= 12'd962;
            12'd778: RELPAGE <= 12'd1484;
            12'd779: RELPAGE <= 12'd2006;
            12'd780: RELPAGE <= 12'd475;
            12'd781: RELPAGE <= 12'd997;
            12'd782: RELPAGE <= 12'd1519;
            12'd783: RELPAGE <= 12'd2041;
            12'd784: RELPAGE <= 12'd510;
            12'd785: RELPAGE <= 12'd1032;
            12'd786: RELPAGE <= 12'd1554;
            12'd787: RELPAGE <= 12'd23;
            12'd788: RELPAGE <= 12'd545;
            12'd789: RELPAGE <= 12'd1067;
            12'd790: RELPAGE <= 12'd1589;
            12'd791: RELPAGE <= 12'd58;
            12'd792: RELPAGE <= 12'd580;
            12'd793: RELPAGE <= 12'd1102;
            12'd794: RELPAGE <= 12'd1624;
            12'd795: RELPAGE <= 12'd93;
            12'd796: RELPAGE <= 12'd615;
            12'd797: RELPAGE <= 12'd1137;
            12'd798: RELPAGE <= 12'd1659;
            12'd799: RELPAGE <= 12'd128;
            12'd800: RELPAGE <= 12'd650;
            12'd801: RELPAGE <= 12'd1172;
            12'd802: RELPAGE <= 12'd1694;
            12'd803: RELPAGE <= 12'd163;
            12'd804: RELPAGE <= 12'd685;
            12'd805: RELPAGE <= 12'd1207;
            12'd806: RELPAGE <= 12'd1729;
            12'd807: RELPAGE <= 12'd198;
            12'd808: RELPAGE <= 12'd720;
            12'd809: RELPAGE <= 12'd1242;
            12'd810: RELPAGE <= 12'd1764;
            12'd811: RELPAGE <= 12'd233;
            12'd812: RELPAGE <= 12'd755;
            12'd813: RELPAGE <= 12'd1277;
            12'd814: RELPAGE <= 12'd1799;
            12'd815: RELPAGE <= 12'd268;
            12'd816: RELPAGE <= 12'd790;
            12'd817: RELPAGE <= 12'd1312;
            12'd818: RELPAGE <= 12'd1834;
            12'd819: RELPAGE <= 12'd303;
            12'd820: RELPAGE <= 12'd825;
            12'd821: RELPAGE <= 12'd1347;
            12'd822: RELPAGE <= 12'd1869;
            12'd823: RELPAGE <= 12'd338;
            12'd824: RELPAGE <= 12'd860;
            12'd825: RELPAGE <= 12'd1382;
            12'd826: RELPAGE <= 12'd1904;
            12'd827: RELPAGE <= 12'd373;
            12'd828: RELPAGE <= 12'd895;
            12'd829: RELPAGE <= 12'd1417;
            12'd830: RELPAGE <= 12'd1939;
            12'd831: RELPAGE <= 12'd408;
            12'd832: RELPAGE <= 12'd930;
            12'd833: RELPAGE <= 12'd1452;
            12'd834: RELPAGE <= 12'd1974;
            12'd835: RELPAGE <= 12'd443;
            12'd836: RELPAGE <= 12'd965;
            12'd837: RELPAGE <= 12'd1487;
            12'd838: RELPAGE <= 12'd2009;
            12'd839: RELPAGE <= 12'd478;
            12'd840: RELPAGE <= 12'd1000;
            12'd841: RELPAGE <= 12'd1522;
            12'd842: RELPAGE <= 12'd2044;
            12'd843: RELPAGE <= 12'd513;
            12'd844: RELPAGE <= 12'd1035;
            12'd845: RELPAGE <= 12'd1557;
            12'd846: RELPAGE <= 12'd26;
            12'd847: RELPAGE <= 12'd548;
            12'd848: RELPAGE <= 12'd1070;
            12'd849: RELPAGE <= 12'd1592;
            12'd850: RELPAGE <= 12'd61;
            12'd851: RELPAGE <= 12'd583;
            12'd852: RELPAGE <= 12'd1105;
            12'd853: RELPAGE <= 12'd1627;
            12'd854: RELPAGE <= 12'd96;
            12'd855: RELPAGE <= 12'd618;
            12'd856: RELPAGE <= 12'd1140;
            12'd857: RELPAGE <= 12'd1662;
            12'd858: RELPAGE <= 12'd131;
            12'd859: RELPAGE <= 12'd653;
            12'd860: RELPAGE <= 12'd1175;
            12'd861: RELPAGE <= 12'd1697;
            12'd862: RELPAGE <= 12'd166;
            12'd863: RELPAGE <= 12'd688;
            12'd864: RELPAGE <= 12'd1210;
            12'd865: RELPAGE <= 12'd1732;
            12'd866: RELPAGE <= 12'd201;
            12'd867: RELPAGE <= 12'd723;
            12'd868: RELPAGE <= 12'd1245;
            12'd869: RELPAGE <= 12'd1767;
            12'd870: RELPAGE <= 12'd236;
            12'd871: RELPAGE <= 12'd758;
            12'd872: RELPAGE <= 12'd1280;
            12'd873: RELPAGE <= 12'd1802;
            12'd874: RELPAGE <= 12'd271;
            12'd875: RELPAGE <= 12'd793;
            12'd876: RELPAGE <= 12'd1315;
            12'd877: RELPAGE <= 12'd1837;
            12'd878: RELPAGE <= 12'd306;
            12'd879: RELPAGE <= 12'd828;
            12'd880: RELPAGE <= 12'd1350;
            12'd881: RELPAGE <= 12'd1872;
            12'd882: RELPAGE <= 12'd341;
            12'd883: RELPAGE <= 12'd863;
            12'd884: RELPAGE <= 12'd1385;
            12'd885: RELPAGE <= 12'd1907;
            12'd886: RELPAGE <= 12'd376;
            12'd887: RELPAGE <= 12'd898;
            12'd888: RELPAGE <= 12'd1420;
            12'd889: RELPAGE <= 12'd1942;
            12'd890: RELPAGE <= 12'd411;
            12'd891: RELPAGE <= 12'd933;
            12'd892: RELPAGE <= 12'd1455;
            12'd893: RELPAGE <= 12'd1977;
            12'd894: RELPAGE <= 12'd446;
            12'd895: RELPAGE <= 12'd968;
            12'd896: RELPAGE <= 12'd1490;
            12'd897: RELPAGE <= 12'd2012;
            12'd898: RELPAGE <= 12'd481;
            12'd899: RELPAGE <= 12'd1003;
            12'd900: RELPAGE <= 12'd1525;
            12'd901: RELPAGE <= 12'd2047;
            12'd902: RELPAGE <= 12'd516;
            12'd903: RELPAGE <= 12'd1038;
            12'd904: RELPAGE <= 12'd1560;
            12'd905: RELPAGE <= 12'd29;
            12'd906: RELPAGE <= 12'd551;
            12'd907: RELPAGE <= 12'd1073;
            12'd908: RELPAGE <= 12'd1595;
            12'd909: RELPAGE <= 12'd64;
            12'd910: RELPAGE <= 12'd586;
            12'd911: RELPAGE <= 12'd1108;
            12'd912: RELPAGE <= 12'd1630;
            12'd913: RELPAGE <= 12'd99;
            12'd914: RELPAGE <= 12'd621;
            12'd915: RELPAGE <= 12'd1143;
            12'd916: RELPAGE <= 12'd1665;
            12'd917: RELPAGE <= 12'd134;
            12'd918: RELPAGE <= 12'd656;
            12'd919: RELPAGE <= 12'd1178;
            12'd920: RELPAGE <= 12'd1700;
            12'd921: RELPAGE <= 12'd169;
            12'd922: RELPAGE <= 12'd691;
            12'd923: RELPAGE <= 12'd1213;
            12'd924: RELPAGE <= 12'd1735;
            12'd925: RELPAGE <= 12'd204;
            12'd926: RELPAGE <= 12'd726;
            12'd927: RELPAGE <= 12'd1248;
            12'd928: RELPAGE <= 12'd1770;
            12'd929: RELPAGE <= 12'd239;
            12'd930: RELPAGE <= 12'd761;
            12'd931: RELPAGE <= 12'd1283;
            12'd932: RELPAGE <= 12'd1805;
            12'd933: RELPAGE <= 12'd274;
            12'd934: RELPAGE <= 12'd796;
            12'd935: RELPAGE <= 12'd1318;
            12'd936: RELPAGE <= 12'd1840;
            12'd937: RELPAGE <= 12'd309;
            12'd938: RELPAGE <= 12'd831;
            12'd939: RELPAGE <= 12'd1353;
            12'd940: RELPAGE <= 12'd1875;
            12'd941: RELPAGE <= 12'd344;
            12'd942: RELPAGE <= 12'd866;
            12'd943: RELPAGE <= 12'd1388;
            12'd944: RELPAGE <= 12'd1910;
            12'd945: RELPAGE <= 12'd379;
            12'd946: RELPAGE <= 12'd901;
            12'd947: RELPAGE <= 12'd1423;
            12'd948: RELPAGE <= 12'd1945;
            12'd949: RELPAGE <= 12'd414;
            12'd950: RELPAGE <= 12'd936;
            12'd951: RELPAGE <= 12'd1458;
            12'd952: RELPAGE <= 12'd1980;
            12'd953: RELPAGE <= 12'd449;
            12'd954: RELPAGE <= 12'd971;
            12'd955: RELPAGE <= 12'd1493;
            12'd956: RELPAGE <= 12'd2015;
            12'd957: RELPAGE <= 12'd484;
            12'd958: RELPAGE <= 12'd1006;
            12'd959: RELPAGE <= 12'd1528;
            12'd960: RELPAGE <= 12'd2050;
            12'd961: RELPAGE <= 12'd519;
            12'd962: RELPAGE <= 12'd1041;
            12'd963: RELPAGE <= 12'd1563;
            12'd964: RELPAGE <= 12'd32;
            12'd965: RELPAGE <= 12'd554;
            12'd966: RELPAGE <= 12'd1076;
            12'd967: RELPAGE <= 12'd1598;
            12'd968: RELPAGE <= 12'd67;
            12'd969: RELPAGE <= 12'd589;
            12'd970: RELPAGE <= 12'd1111;
            12'd971: RELPAGE <= 12'd1633;
            12'd972: RELPAGE <= 12'd102;
            12'd973: RELPAGE <= 12'd624;
            12'd974: RELPAGE <= 12'd1146;
            12'd975: RELPAGE <= 12'd1668;
            12'd976: RELPAGE <= 12'd137;
            12'd977: RELPAGE <= 12'd659;
            12'd978: RELPAGE <= 12'd1181;
            12'd979: RELPAGE <= 12'd1703;
            12'd980: RELPAGE <= 12'd172;
            12'd981: RELPAGE <= 12'd694;
            12'd982: RELPAGE <= 12'd1216;
            12'd983: RELPAGE <= 12'd1738;
            12'd984: RELPAGE <= 12'd207;
            12'd985: RELPAGE <= 12'd729;
            12'd986: RELPAGE <= 12'd1251;
            12'd987: RELPAGE <= 12'd1773;
            12'd988: RELPAGE <= 12'd242;
            12'd989: RELPAGE <= 12'd764;
            12'd990: RELPAGE <= 12'd1286;
            12'd991: RELPAGE <= 12'd1808;
            12'd992: RELPAGE <= 12'd277;
            12'd993: RELPAGE <= 12'd799;
            12'd994: RELPAGE <= 12'd1321;
            12'd995: RELPAGE <= 12'd1843;
            12'd996: RELPAGE <= 12'd312;
            12'd997: RELPAGE <= 12'd834;
            12'd998: RELPAGE <= 12'd1356;
            12'd999: RELPAGE <= 12'd1878;
            12'd1000: RELPAGE <= 12'd347;
            12'd1001: RELPAGE <= 12'd869;
            12'd1002: RELPAGE <= 12'd1391;
            12'd1003: RELPAGE <= 12'd1913;
            12'd1004: RELPAGE <= 12'd382;
            12'd1005: RELPAGE <= 12'd904;
            12'd1006: RELPAGE <= 12'd1426;
            12'd1007: RELPAGE <= 12'd1948;
            12'd1008: RELPAGE <= 12'd417;
            12'd1009: RELPAGE <= 12'd939;
            12'd1010: RELPAGE <= 12'd1461;
            12'd1011: RELPAGE <= 12'd1983;
            12'd1012: RELPAGE <= 12'd452;
            12'd1013: RELPAGE <= 12'd974;
            12'd1014: RELPAGE <= 12'd1496;
            12'd1015: RELPAGE <= 12'd2018;
            12'd1016: RELPAGE <= 12'd487;
            12'd1017: RELPAGE <= 12'd1009;
            12'd1018: RELPAGE <= 12'd1531;
            12'd1019: RELPAGE <= 12'd0;
            12'd1020: RELPAGE <= 12'd522;
            12'd1021: RELPAGE <= 12'd1044;
            12'd1022: RELPAGE <= 12'd1566;
            12'd1023: RELPAGE <= 12'd35;
            12'd1024: RELPAGE <= 12'd557;
            12'd1025: RELPAGE <= 12'd1079;
            12'd1026: RELPAGE <= 12'd1601;
            12'd1027: RELPAGE <= 12'd70;
            12'd1028: RELPAGE <= 12'd592;
            12'd1029: RELPAGE <= 12'd1114;
            12'd1030: RELPAGE <= 12'd1636;
            12'd1031: RELPAGE <= 12'd105;
            12'd1032: RELPAGE <= 12'd627;
            12'd1033: RELPAGE <= 12'd1149;
            12'd1034: RELPAGE <= 12'd1671;
            12'd1035: RELPAGE <= 12'd140;
            12'd1036: RELPAGE <= 12'd662;
            12'd1037: RELPAGE <= 12'd1184;
            12'd1038: RELPAGE <= 12'd1706;
            12'd1039: RELPAGE <= 12'd175;
            12'd1040: RELPAGE <= 12'd697;
            12'd1041: RELPAGE <= 12'd1219;
            12'd1042: RELPAGE <= 12'd1741;
            12'd1043: RELPAGE <= 12'd210;
            12'd1044: RELPAGE <= 12'd732;
            12'd1045: RELPAGE <= 12'd1254;
            12'd1046: RELPAGE <= 12'd1776;
            12'd1047: RELPAGE <= 12'd245;
            12'd1048: RELPAGE <= 12'd767;
            12'd1049: RELPAGE <= 12'd1289;
            12'd1050: RELPAGE <= 12'd1811;
            12'd1051: RELPAGE <= 12'd280;
            12'd1052: RELPAGE <= 12'd802;
            12'd1053: RELPAGE <= 12'd1324;
            12'd1054: RELPAGE <= 12'd1846;
            12'd1055: RELPAGE <= 12'd315;
            12'd1056: RELPAGE <= 12'd837;
            12'd1057: RELPAGE <= 12'd1359;
            12'd1058: RELPAGE <= 12'd1881;
            12'd1059: RELPAGE <= 12'd350;
            12'd1060: RELPAGE <= 12'd872;
            12'd1061: RELPAGE <= 12'd1394;
            12'd1062: RELPAGE <= 12'd1916;
            12'd1063: RELPAGE <= 12'd385;
            12'd1064: RELPAGE <= 12'd907;
            12'd1065: RELPAGE <= 12'd1429;
            12'd1066: RELPAGE <= 12'd1951;
            12'd1067: RELPAGE <= 12'd420;
            12'd1068: RELPAGE <= 12'd942;
            12'd1069: RELPAGE <= 12'd1464;
            12'd1070: RELPAGE <= 12'd1986;
            12'd1071: RELPAGE <= 12'd455;
            12'd1072: RELPAGE <= 12'd977;
            12'd1073: RELPAGE <= 12'd1499;
            12'd1074: RELPAGE <= 12'd2021;
            12'd1075: RELPAGE <= 12'd490;
            12'd1076: RELPAGE <= 12'd1012;
            12'd1077: RELPAGE <= 12'd1534;
            12'd1078: RELPAGE <= 12'd3;
            12'd1079: RELPAGE <= 12'd525;
            12'd1080: RELPAGE <= 12'd1047;
            12'd1081: RELPAGE <= 12'd1569;
            12'd1082: RELPAGE <= 12'd38;
            12'd1083: RELPAGE <= 12'd560;
            12'd1084: RELPAGE <= 12'd1082;
            12'd1085: RELPAGE <= 12'd1604;
            12'd1086: RELPAGE <= 12'd73;
            12'd1087: RELPAGE <= 12'd595;
            12'd1088: RELPAGE <= 12'd1117;
            12'd1089: RELPAGE <= 12'd1639;
            12'd1090: RELPAGE <= 12'd108;
            12'd1091: RELPAGE <= 12'd630;
            12'd1092: RELPAGE <= 12'd1152;
            12'd1093: RELPAGE <= 12'd1674;
            12'd1094: RELPAGE <= 12'd143;
            12'd1095: RELPAGE <= 12'd665;
            12'd1096: RELPAGE <= 12'd1187;
            12'd1097: RELPAGE <= 12'd1709;
            12'd1098: RELPAGE <= 12'd178;
            12'd1099: RELPAGE <= 12'd700;
            12'd1100: RELPAGE <= 12'd1222;
            12'd1101: RELPAGE <= 12'd1744;
            12'd1102: RELPAGE <= 12'd213;
            12'd1103: RELPAGE <= 12'd735;
            12'd1104: RELPAGE <= 12'd1257;
            12'd1105: RELPAGE <= 12'd1779;
            12'd1106: RELPAGE <= 12'd248;
            12'd1107: RELPAGE <= 12'd770;
            12'd1108: RELPAGE <= 12'd1292;
            12'd1109: RELPAGE <= 12'd1814;
            12'd1110: RELPAGE <= 12'd283;
            12'd1111: RELPAGE <= 12'd805;
            12'd1112: RELPAGE <= 12'd1327;
            12'd1113: RELPAGE <= 12'd1849;
            12'd1114: RELPAGE <= 12'd318;
            12'd1115: RELPAGE <= 12'd840;
            12'd1116: RELPAGE <= 12'd1362;
            12'd1117: RELPAGE <= 12'd1884;
            12'd1118: RELPAGE <= 12'd353;
            12'd1119: RELPAGE <= 12'd875;
            12'd1120: RELPAGE <= 12'd1397;
            12'd1121: RELPAGE <= 12'd1919;
            12'd1122: RELPAGE <= 12'd388;
            12'd1123: RELPAGE <= 12'd910;
            12'd1124: RELPAGE <= 12'd1432;
            12'd1125: RELPAGE <= 12'd1954;
            12'd1126: RELPAGE <= 12'd423;
            12'd1127: RELPAGE <= 12'd945;
            12'd1128: RELPAGE <= 12'd1467;
            12'd1129: RELPAGE <= 12'd1989;
            12'd1130: RELPAGE <= 12'd458;
            12'd1131: RELPAGE <= 12'd980;
            12'd1132: RELPAGE <= 12'd1502;
            12'd1133: RELPAGE <= 12'd2024;
            12'd1134: RELPAGE <= 12'd493;
            12'd1135: RELPAGE <= 12'd1015;
            12'd1136: RELPAGE <= 12'd1537;
            12'd1137: RELPAGE <= 12'd6;
            12'd1138: RELPAGE <= 12'd528;
            12'd1139: RELPAGE <= 12'd1050;
            12'd1140: RELPAGE <= 12'd1572;
            12'd1141: RELPAGE <= 12'd41;
            12'd1142: RELPAGE <= 12'd563;
            12'd1143: RELPAGE <= 12'd1085;
            12'd1144: RELPAGE <= 12'd1607;
            12'd1145: RELPAGE <= 12'd76;
            12'd1146: RELPAGE <= 12'd598;
            12'd1147: RELPAGE <= 12'd1120;
            12'd1148: RELPAGE <= 12'd1642;
            12'd1149: RELPAGE <= 12'd111;
            12'd1150: RELPAGE <= 12'd633;
            12'd1151: RELPAGE <= 12'd1155;
            12'd1152: RELPAGE <= 12'd1677;
            12'd1153: RELPAGE <= 12'd146;
            12'd1154: RELPAGE <= 12'd668;
            12'd1155: RELPAGE <= 12'd1190;
            12'd1156: RELPAGE <= 12'd1712;
            12'd1157: RELPAGE <= 12'd181;
            12'd1158: RELPAGE <= 12'd703;
            12'd1159: RELPAGE <= 12'd1225;
            12'd1160: RELPAGE <= 12'd1747;
            12'd1161: RELPAGE <= 12'd216;
            12'd1162: RELPAGE <= 12'd738;
            12'd1163: RELPAGE <= 12'd1260;
            12'd1164: RELPAGE <= 12'd1782;
            12'd1165: RELPAGE <= 12'd251;
            12'd1166: RELPAGE <= 12'd773;
            12'd1167: RELPAGE <= 12'd1295;
            12'd1168: RELPAGE <= 12'd1817;
            12'd1169: RELPAGE <= 12'd286;
            12'd1170: RELPAGE <= 12'd808;
            12'd1171: RELPAGE <= 12'd1330;
            12'd1172: RELPAGE <= 12'd1852;
            12'd1173: RELPAGE <= 12'd321;
            12'd1174: RELPAGE <= 12'd843;
            12'd1175: RELPAGE <= 12'd1365;
            12'd1176: RELPAGE <= 12'd1887;
            12'd1177: RELPAGE <= 12'd356;
            12'd1178: RELPAGE <= 12'd878;
            12'd1179: RELPAGE <= 12'd1400;
            12'd1180: RELPAGE <= 12'd1922;
            12'd1181: RELPAGE <= 12'd391;
            12'd1182: RELPAGE <= 12'd913;
            12'd1183: RELPAGE <= 12'd1435;
            12'd1184: RELPAGE <= 12'd1957;
            12'd1185: RELPAGE <= 12'd426;
            12'd1186: RELPAGE <= 12'd948;
            12'd1187: RELPAGE <= 12'd1470;
            12'd1188: RELPAGE <= 12'd1992;
            12'd1189: RELPAGE <= 12'd461;
            12'd1190: RELPAGE <= 12'd983;
            12'd1191: RELPAGE <= 12'd1505;
            12'd1192: RELPAGE <= 12'd2027;
            12'd1193: RELPAGE <= 12'd496;
            12'd1194: RELPAGE <= 12'd1018;
            12'd1195: RELPAGE <= 12'd1540;
            12'd1196: RELPAGE <= 12'd9;
            12'd1197: RELPAGE <= 12'd531;
            12'd1198: RELPAGE <= 12'd1053;
            12'd1199: RELPAGE <= 12'd1575;
            12'd1200: RELPAGE <= 12'd44;
            12'd1201: RELPAGE <= 12'd566;
            12'd1202: RELPAGE <= 12'd1088;
            12'd1203: RELPAGE <= 12'd1610;
            12'd1204: RELPAGE <= 12'd79;
            12'd1205: RELPAGE <= 12'd601;
            12'd1206: RELPAGE <= 12'd1123;
            12'd1207: RELPAGE <= 12'd1645;
            12'd1208: RELPAGE <= 12'd114;
            12'd1209: RELPAGE <= 12'd636;
            12'd1210: RELPAGE <= 12'd1158;
            12'd1211: RELPAGE <= 12'd1680;
            12'd1212: RELPAGE <= 12'd149;
            12'd1213: RELPAGE <= 12'd671;
            12'd1214: RELPAGE <= 12'd1193;
            12'd1215: RELPAGE <= 12'd1715;
            12'd1216: RELPAGE <= 12'd184;
            12'd1217: RELPAGE <= 12'd706;
            12'd1218: RELPAGE <= 12'd1228;
            12'd1219: RELPAGE <= 12'd1750;
            12'd1220: RELPAGE <= 12'd219;
            12'd1221: RELPAGE <= 12'd741;
            12'd1222: RELPAGE <= 12'd1263;
            12'd1223: RELPAGE <= 12'd1785;
            12'd1224: RELPAGE <= 12'd254;
            12'd1225: RELPAGE <= 12'd776;
            12'd1226: RELPAGE <= 12'd1298;
            12'd1227: RELPAGE <= 12'd1820;
            12'd1228: RELPAGE <= 12'd289;
            12'd1229: RELPAGE <= 12'd811;
            12'd1230: RELPAGE <= 12'd1333;
            12'd1231: RELPAGE <= 12'd1855;
            12'd1232: RELPAGE <= 12'd324;
            12'd1233: RELPAGE <= 12'd846;
            12'd1234: RELPAGE <= 12'd1368;
            12'd1235: RELPAGE <= 12'd1890;
            12'd1236: RELPAGE <= 12'd359;
            12'd1237: RELPAGE <= 12'd881;
            12'd1238: RELPAGE <= 12'd1403;
            12'd1239: RELPAGE <= 12'd1925;
            12'd1240: RELPAGE <= 12'd394;
            12'd1241: RELPAGE <= 12'd916;
            12'd1242: RELPAGE <= 12'd1438;
            12'd1243: RELPAGE <= 12'd1960;
            12'd1244: RELPAGE <= 12'd429;
            12'd1245: RELPAGE <= 12'd951;
            12'd1246: RELPAGE <= 12'd1473;
            12'd1247: RELPAGE <= 12'd1995;
            12'd1248: RELPAGE <= 12'd464;
            12'd1249: RELPAGE <= 12'd986;
            12'd1250: RELPAGE <= 12'd1508;
            12'd1251: RELPAGE <= 12'd2030;
            12'd1252: RELPAGE <= 12'd499;
            12'd1253: RELPAGE <= 12'd1021;
            12'd1254: RELPAGE <= 12'd1543;
            12'd1255: RELPAGE <= 12'd12;
            12'd1256: RELPAGE <= 12'd534;
            12'd1257: RELPAGE <= 12'd1056;
            12'd1258: RELPAGE <= 12'd1578;
            12'd1259: RELPAGE <= 12'd47;
            12'd1260: RELPAGE <= 12'd569;
            12'd1261: RELPAGE <= 12'd1091;
            12'd1262: RELPAGE <= 12'd1613;
            12'd1263: RELPAGE <= 12'd82;
            12'd1264: RELPAGE <= 12'd604;
            12'd1265: RELPAGE <= 12'd1126;
            12'd1266: RELPAGE <= 12'd1648;
            12'd1267: RELPAGE <= 12'd117;
            12'd1268: RELPAGE <= 12'd639;
            12'd1269: RELPAGE <= 12'd1161;
            12'd1270: RELPAGE <= 12'd1683;
            12'd1271: RELPAGE <= 12'd152;
            12'd1272: RELPAGE <= 12'd674;
            12'd1273: RELPAGE <= 12'd1196;
            12'd1274: RELPAGE <= 12'd1718;
            12'd1275: RELPAGE <= 12'd187;
            12'd1276: RELPAGE <= 12'd709;
            12'd1277: RELPAGE <= 12'd1231;
            12'd1278: RELPAGE <= 12'd1753;
            12'd1279: RELPAGE <= 12'd222;
            12'd1280: RELPAGE <= 12'd744;
            12'd1281: RELPAGE <= 12'd1266;
            12'd1282: RELPAGE <= 12'd1788;
            12'd1283: RELPAGE <= 12'd257;
            12'd1284: RELPAGE <= 12'd779;
            12'd1285: RELPAGE <= 12'd1301;
            12'd1286: RELPAGE <= 12'd1823;
            12'd1287: RELPAGE <= 12'd292;
            12'd1288: RELPAGE <= 12'd814;
            12'd1289: RELPAGE <= 12'd1336;
            12'd1290: RELPAGE <= 12'd1858;
            12'd1291: RELPAGE <= 12'd327;
            12'd1292: RELPAGE <= 12'd849;
            12'd1293: RELPAGE <= 12'd1371;
            12'd1294: RELPAGE <= 12'd1893;
            12'd1295: RELPAGE <= 12'd362;
            12'd1296: RELPAGE <= 12'd884;
            12'd1297: RELPAGE <= 12'd1406;
            12'd1298: RELPAGE <= 12'd1928;
            12'd1299: RELPAGE <= 12'd397;
            12'd1300: RELPAGE <= 12'd919;
            12'd1301: RELPAGE <= 12'd1441;
            12'd1302: RELPAGE <= 12'd1963;
            12'd1303: RELPAGE <= 12'd432;
            12'd1304: RELPAGE <= 12'd954;
            12'd1305: RELPAGE <= 12'd1476;
            12'd1306: RELPAGE <= 12'd1998;
            12'd1307: RELPAGE <= 12'd467;
            12'd1308: RELPAGE <= 12'd989;
            12'd1309: RELPAGE <= 12'd1511;
            12'd1310: RELPAGE <= 12'd2033;
            12'd1311: RELPAGE <= 12'd502;
            12'd1312: RELPAGE <= 12'd1024;
            12'd1313: RELPAGE <= 12'd1546;
            12'd1314: RELPAGE <= 12'd15;
            12'd1315: RELPAGE <= 12'd537;
            12'd1316: RELPAGE <= 12'd1059;
            12'd1317: RELPAGE <= 12'd1581;
            12'd1318: RELPAGE <= 12'd50;
            12'd1319: RELPAGE <= 12'd572;
            12'd1320: RELPAGE <= 12'd1094;
            12'd1321: RELPAGE <= 12'd1616;
            12'd1322: RELPAGE <= 12'd85;
            12'd1323: RELPAGE <= 12'd607;
            12'd1324: RELPAGE <= 12'd1129;
            12'd1325: RELPAGE <= 12'd1651;
            12'd1326: RELPAGE <= 12'd120;
            12'd1327: RELPAGE <= 12'd642;
            12'd1328: RELPAGE <= 12'd1164;
            12'd1329: RELPAGE <= 12'd1686;
            12'd1330: RELPAGE <= 12'd155;
            12'd1331: RELPAGE <= 12'd677;
            12'd1332: RELPAGE <= 12'd1199;
            12'd1333: RELPAGE <= 12'd1721;
            12'd1334: RELPAGE <= 12'd190;
            12'd1335: RELPAGE <= 12'd712;
            12'd1336: RELPAGE <= 12'd1234;
            12'd1337: RELPAGE <= 12'd1756;
            12'd1338: RELPAGE <= 12'd225;
            12'd1339: RELPAGE <= 12'd747;
            12'd1340: RELPAGE <= 12'd1269;
            12'd1341: RELPAGE <= 12'd1791;
            12'd1342: RELPAGE <= 12'd260;
            12'd1343: RELPAGE <= 12'd782;
            12'd1344: RELPAGE <= 12'd1304;
            12'd1345: RELPAGE <= 12'd1826;
            12'd1346: RELPAGE <= 12'd295;
            12'd1347: RELPAGE <= 12'd817;
            12'd1348: RELPAGE <= 12'd1339;
            12'd1349: RELPAGE <= 12'd1861;
            12'd1350: RELPAGE <= 12'd330;
            12'd1351: RELPAGE <= 12'd852;
            12'd1352: RELPAGE <= 12'd1374;
            12'd1353: RELPAGE <= 12'd1896;
            12'd1354: RELPAGE <= 12'd365;
            12'd1355: RELPAGE <= 12'd887;
            12'd1356: RELPAGE <= 12'd1409;
            12'd1357: RELPAGE <= 12'd1931;
            12'd1358: RELPAGE <= 12'd400;
            12'd1359: RELPAGE <= 12'd922;
            12'd1360: RELPAGE <= 12'd1444;
            12'd1361: RELPAGE <= 12'd1966;
            12'd1362: RELPAGE <= 12'd435;
            12'd1363: RELPAGE <= 12'd957;
            12'd1364: RELPAGE <= 12'd1479;
            12'd1365: RELPAGE <= 12'd2001;
            12'd1366: RELPAGE <= 12'd470;
            12'd1367: RELPAGE <= 12'd992;
            12'd1368: RELPAGE <= 12'd1514;
            12'd1369: RELPAGE <= 12'd2036;
            12'd1370: RELPAGE <= 12'd505;
            12'd1371: RELPAGE <= 12'd1027;
            12'd1372: RELPAGE <= 12'd1549;
            12'd1373: RELPAGE <= 12'd18;
            12'd1374: RELPAGE <= 12'd540;
            12'd1375: RELPAGE <= 12'd1062;
            12'd1376: RELPAGE <= 12'd1584;
            12'd1377: RELPAGE <= 12'd53;
            12'd1378: RELPAGE <= 12'd575;
            12'd1379: RELPAGE <= 12'd1097;
            12'd1380: RELPAGE <= 12'd1619;
            12'd1381: RELPAGE <= 12'd88;
            12'd1382: RELPAGE <= 12'd610;
            12'd1383: RELPAGE <= 12'd1132;
            12'd1384: RELPAGE <= 12'd1654;
            12'd1385: RELPAGE <= 12'd123;
            12'd1386: RELPAGE <= 12'd645;
            12'd1387: RELPAGE <= 12'd1167;
            12'd1388: RELPAGE <= 12'd1689;
            12'd1389: RELPAGE <= 12'd158;
            12'd1390: RELPAGE <= 12'd680;
            12'd1391: RELPAGE <= 12'd1202;
            12'd1392: RELPAGE <= 12'd1724;
            12'd1393: RELPAGE <= 12'd193;
            12'd1394: RELPAGE <= 12'd715;
            12'd1395: RELPAGE <= 12'd1237;
            12'd1396: RELPAGE <= 12'd1759;
            12'd1397: RELPAGE <= 12'd228;
            12'd1398: RELPAGE <= 12'd750;
            12'd1399: RELPAGE <= 12'd1272;
            12'd1400: RELPAGE <= 12'd1794;
            12'd1401: RELPAGE <= 12'd263;
            12'd1402: RELPAGE <= 12'd785;
            12'd1403: RELPAGE <= 12'd1307;
            12'd1404: RELPAGE <= 12'd1829;
            12'd1405: RELPAGE <= 12'd298;
            12'd1406: RELPAGE <= 12'd820;
            12'd1407: RELPAGE <= 12'd1342;
            12'd1408: RELPAGE <= 12'd1864;
            12'd1409: RELPAGE <= 12'd333;
            12'd1410: RELPAGE <= 12'd855;
            12'd1411: RELPAGE <= 12'd1377;
            12'd1412: RELPAGE <= 12'd1899;
            12'd1413: RELPAGE <= 12'd368;
            12'd1414: RELPAGE <= 12'd890;
            12'd1415: RELPAGE <= 12'd1412;
            12'd1416: RELPAGE <= 12'd1934;
            12'd1417: RELPAGE <= 12'd403;
            12'd1418: RELPAGE <= 12'd925;
            12'd1419: RELPAGE <= 12'd1447;
            12'd1420: RELPAGE <= 12'd1969;
            12'd1421: RELPAGE <= 12'd438;
            12'd1422: RELPAGE <= 12'd960;
            12'd1423: RELPAGE <= 12'd1482;
            12'd1424: RELPAGE <= 12'd2004;
            12'd1425: RELPAGE <= 12'd473;
            12'd1426: RELPAGE <= 12'd995;
            12'd1427: RELPAGE <= 12'd1517;
            12'd1428: RELPAGE <= 12'd2039;
            12'd1429: RELPAGE <= 12'd508;
            12'd1430: RELPAGE <= 12'd1030;
            12'd1431: RELPAGE <= 12'd1552;
            12'd1432: RELPAGE <= 12'd21;
            12'd1433: RELPAGE <= 12'd543;
            12'd1434: RELPAGE <= 12'd1065;
            12'd1435: RELPAGE <= 12'd1587;
            12'd1436: RELPAGE <= 12'd56;
            12'd1437: RELPAGE <= 12'd578;
            12'd1438: RELPAGE <= 12'd1100;
            12'd1439: RELPAGE <= 12'd1622;
            12'd1440: RELPAGE <= 12'd91;
            12'd1441: RELPAGE <= 12'd613;
            12'd1442: RELPAGE <= 12'd1135;
            12'd1443: RELPAGE <= 12'd1657;
            12'd1444: RELPAGE <= 12'd126;
            12'd1445: RELPAGE <= 12'd648;
            12'd1446: RELPAGE <= 12'd1170;
            12'd1447: RELPAGE <= 12'd1692;
            12'd1448: RELPAGE <= 12'd161;
            12'd1449: RELPAGE <= 12'd683;
            12'd1450: RELPAGE <= 12'd1205;
            12'd1451: RELPAGE <= 12'd1727;
            12'd1452: RELPAGE <= 12'd196;
            12'd1453: RELPAGE <= 12'd718;
            12'd1454: RELPAGE <= 12'd1240;
            12'd1455: RELPAGE <= 12'd1762;
            12'd1456: RELPAGE <= 12'd231;
            12'd1457: RELPAGE <= 12'd753;
            12'd1458: RELPAGE <= 12'd1275;
            12'd1459: RELPAGE <= 12'd1797;
            12'd1460: RELPAGE <= 12'd266;
            12'd1461: RELPAGE <= 12'd788;
            12'd1462: RELPAGE <= 12'd1310;
            12'd1463: RELPAGE <= 12'd1832;
            12'd1464: RELPAGE <= 12'd301;
            12'd1465: RELPAGE <= 12'd823;
            12'd1466: RELPAGE <= 12'd1345;
            12'd1467: RELPAGE <= 12'd1867;
            12'd1468: RELPAGE <= 12'd336;
            12'd1469: RELPAGE <= 12'd858;
            12'd1470: RELPAGE <= 12'd1380;
            12'd1471: RELPAGE <= 12'd1902;
            12'd1472: RELPAGE <= 12'd371;
            12'd1473: RELPAGE <= 12'd893;
            12'd1474: RELPAGE <= 12'd1415;
            12'd1475: RELPAGE <= 12'd1937;
            12'd1476: RELPAGE <= 12'd406;
            12'd1477: RELPAGE <= 12'd928;
            12'd1478: RELPAGE <= 12'd1450;
            12'd1479: RELPAGE <= 12'd1972;
            12'd1480: RELPAGE <= 12'd441;
            12'd1481: RELPAGE <= 12'd963;
            12'd1482: RELPAGE <= 12'd1485;
            12'd1483: RELPAGE <= 12'd2007;
            12'd1484: RELPAGE <= 12'd476;
            12'd1485: RELPAGE <= 12'd998;
            12'd1486: RELPAGE <= 12'd1520;
            12'd1487: RELPAGE <= 12'd2042;
            12'd1488: RELPAGE <= 12'd511;
            12'd1489: RELPAGE <= 12'd1033;
            12'd1490: RELPAGE <= 12'd1555;
            12'd1491: RELPAGE <= 12'd24;
            12'd1492: RELPAGE <= 12'd546;
            12'd1493: RELPAGE <= 12'd1068;
            12'd1494: RELPAGE <= 12'd1590;
            12'd1495: RELPAGE <= 12'd59;
            12'd1496: RELPAGE <= 12'd581;
            12'd1497: RELPAGE <= 12'd1103;
            12'd1498: RELPAGE <= 12'd1625;
            12'd1499: RELPAGE <= 12'd94;
            12'd1500: RELPAGE <= 12'd616;
            12'd1501: RELPAGE <= 12'd1138;
            12'd1502: RELPAGE <= 12'd1660;
            12'd1503: RELPAGE <= 12'd129;
            12'd1504: RELPAGE <= 12'd651;
            12'd1505: RELPAGE <= 12'd1173;
            12'd1506: RELPAGE <= 12'd1695;
            12'd1507: RELPAGE <= 12'd164;
            12'd1508: RELPAGE <= 12'd686;
            12'd1509: RELPAGE <= 12'd1208;
            12'd1510: RELPAGE <= 12'd1730;
            12'd1511: RELPAGE <= 12'd199;
            12'd1512: RELPAGE <= 12'd721;
            12'd1513: RELPAGE <= 12'd1243;
            12'd1514: RELPAGE <= 12'd1765;
            12'd1515: RELPAGE <= 12'd234;
            12'd1516: RELPAGE <= 12'd756;
            12'd1517: RELPAGE <= 12'd1278;
            12'd1518: RELPAGE <= 12'd1800;
            12'd1519: RELPAGE <= 12'd269;
            12'd1520: RELPAGE <= 12'd791;
            12'd1521: RELPAGE <= 12'd1313;
            12'd1522: RELPAGE <= 12'd1835;
            12'd1523: RELPAGE <= 12'd304;
            12'd1524: RELPAGE <= 12'd826;
            12'd1525: RELPAGE <= 12'd1348;
            12'd1526: RELPAGE <= 12'd1870;
            12'd1527: RELPAGE <= 12'd339;
            12'd1528: RELPAGE <= 12'd861;
            12'd1529: RELPAGE <= 12'd1383;
            12'd1530: RELPAGE <= 12'd1905;
            12'd1531: RELPAGE <= 12'd374;
            12'd1532: RELPAGE <= 12'd896;
            12'd1533: RELPAGE <= 12'd1418;
            12'd1534: RELPAGE <= 12'd1940;
            12'd1535: RELPAGE <= 12'd409;
            12'd1536: RELPAGE <= 12'd931;
            12'd1537: RELPAGE <= 12'd1453;
            12'd1538: RELPAGE <= 12'd1975;
            12'd1539: RELPAGE <= 12'd444;
            12'd1540: RELPAGE <= 12'd966;
            12'd1541: RELPAGE <= 12'd1488;
            12'd1542: RELPAGE <= 12'd2010;
            12'd1543: RELPAGE <= 12'd479;
            12'd1544: RELPAGE <= 12'd1001;
            12'd1545: RELPAGE <= 12'd1523;
            12'd1546: RELPAGE <= 12'd2045;
            12'd1547: RELPAGE <= 12'd514;
            12'd1548: RELPAGE <= 12'd1036;
            12'd1549: RELPAGE <= 12'd1558;
            12'd1550: RELPAGE <= 12'd27;
            12'd1551: RELPAGE <= 12'd549;
            12'd1552: RELPAGE <= 12'd1071;
            12'd1553: RELPAGE <= 12'd1593;
            12'd1554: RELPAGE <= 12'd62;
            12'd1555: RELPAGE <= 12'd584;
            12'd1556: RELPAGE <= 12'd1106;
            12'd1557: RELPAGE <= 12'd1628;
            12'd1558: RELPAGE <= 12'd97;
            12'd1559: RELPAGE <= 12'd619;
            12'd1560: RELPAGE <= 12'd1141;
            12'd1561: RELPAGE <= 12'd1663;
            12'd1562: RELPAGE <= 12'd132;
            12'd1563: RELPAGE <= 12'd654;
            12'd1564: RELPAGE <= 12'd1176;
            12'd1565: RELPAGE <= 12'd1698;
            12'd1566: RELPAGE <= 12'd167;
            12'd1567: RELPAGE <= 12'd689;
            12'd1568: RELPAGE <= 12'd1211;
            12'd1569: RELPAGE <= 12'd1733;
            12'd1570: RELPAGE <= 12'd202;
            12'd1571: RELPAGE <= 12'd724;
            12'd1572: RELPAGE <= 12'd1246;
            12'd1573: RELPAGE <= 12'd1768;
            12'd1574: RELPAGE <= 12'd237;
            12'd1575: RELPAGE <= 12'd759;
            12'd1576: RELPAGE <= 12'd1281;
            12'd1577: RELPAGE <= 12'd1803;
            12'd1578: RELPAGE <= 12'd272;
            12'd1579: RELPAGE <= 12'd794;
            12'd1580: RELPAGE <= 12'd1316;
            12'd1581: RELPAGE <= 12'd1838;
            12'd1582: RELPAGE <= 12'd307;
            12'd1583: RELPAGE <= 12'd829;
            12'd1584: RELPAGE <= 12'd1351;
            12'd1585: RELPAGE <= 12'd1873;
            12'd1586: RELPAGE <= 12'd342;
            12'd1587: RELPAGE <= 12'd864;
            12'd1588: RELPAGE <= 12'd1386;
            12'd1589: RELPAGE <= 12'd1908;
            12'd1590: RELPAGE <= 12'd377;
            12'd1591: RELPAGE <= 12'd899;
            12'd1592: RELPAGE <= 12'd1421;
            12'd1593: RELPAGE <= 12'd1943;
            12'd1594: RELPAGE <= 12'd412;
            12'd1595: RELPAGE <= 12'd934;
            12'd1596: RELPAGE <= 12'd1456;
            12'd1597: RELPAGE <= 12'd1978;
            12'd1598: RELPAGE <= 12'd447;
            12'd1599: RELPAGE <= 12'd969;
            12'd1600: RELPAGE <= 12'd1491;
            12'd1601: RELPAGE <= 12'd2013;
            12'd1602: RELPAGE <= 12'd482;
            12'd1603: RELPAGE <= 12'd1004;
            12'd1604: RELPAGE <= 12'd1526;
            12'd1605: RELPAGE <= 12'd2048;
            12'd1606: RELPAGE <= 12'd517;
            12'd1607: RELPAGE <= 12'd1039;
            12'd1608: RELPAGE <= 12'd1561;
            12'd1609: RELPAGE <= 12'd30;
            12'd1610: RELPAGE <= 12'd552;
            12'd1611: RELPAGE <= 12'd1074;
            12'd1612: RELPAGE <= 12'd1596;
            12'd1613: RELPAGE <= 12'd65;
            12'd1614: RELPAGE <= 12'd587;
            12'd1615: RELPAGE <= 12'd1109;
            12'd1616: RELPAGE <= 12'd1631;
            12'd1617: RELPAGE <= 12'd100;
            12'd1618: RELPAGE <= 12'd622;
            12'd1619: RELPAGE <= 12'd1144;
            12'd1620: RELPAGE <= 12'd1666;
            12'd1621: RELPAGE <= 12'd135;
            12'd1622: RELPAGE <= 12'd657;
            12'd1623: RELPAGE <= 12'd1179;
            12'd1624: RELPAGE <= 12'd1701;
            12'd1625: RELPAGE <= 12'd170;
            12'd1626: RELPAGE <= 12'd692;
            12'd1627: RELPAGE <= 12'd1214;
            12'd1628: RELPAGE <= 12'd1736;
            12'd1629: RELPAGE <= 12'd205;
            12'd1630: RELPAGE <= 12'd727;
            12'd1631: RELPAGE <= 12'd1249;
            12'd1632: RELPAGE <= 12'd1771;
            12'd1633: RELPAGE <= 12'd240;
            12'd1634: RELPAGE <= 12'd762;
            12'd1635: RELPAGE <= 12'd1284;
            12'd1636: RELPAGE <= 12'd1806;
            12'd1637: RELPAGE <= 12'd275;
            12'd1638: RELPAGE <= 12'd797;
            12'd1639: RELPAGE <= 12'd1319;
            12'd1640: RELPAGE <= 12'd1841;
            12'd1641: RELPAGE <= 12'd310;
            12'd1642: RELPAGE <= 12'd832;
            12'd1643: RELPAGE <= 12'd1354;
            12'd1644: RELPAGE <= 12'd1876;
            12'd1645: RELPAGE <= 12'd345;
            12'd1646: RELPAGE <= 12'd867;
            12'd1647: RELPAGE <= 12'd1389;
            12'd1648: RELPAGE <= 12'd1911;
            12'd1649: RELPAGE <= 12'd380;
            12'd1650: RELPAGE <= 12'd902;
            12'd1651: RELPAGE <= 12'd1424;
            12'd1652: RELPAGE <= 12'd1946;
            12'd1653: RELPAGE <= 12'd415;
            12'd1654: RELPAGE <= 12'd937;
            12'd1655: RELPAGE <= 12'd1459;
            12'd1656: RELPAGE <= 12'd1981;
            12'd1657: RELPAGE <= 12'd450;
            12'd1658: RELPAGE <= 12'd972;
            12'd1659: RELPAGE <= 12'd1494;
            12'd1660: RELPAGE <= 12'd2016;
            12'd1661: RELPAGE <= 12'd485;
            12'd1662: RELPAGE <= 12'd1007;
            12'd1663: RELPAGE <= 12'd1529;
            12'd1664: RELPAGE <= 12'd2051;
            12'd1665: RELPAGE <= 12'd520;
            12'd1666: RELPAGE <= 12'd1042;
            12'd1667: RELPAGE <= 12'd1564;
            12'd1668: RELPAGE <= 12'd33;
            12'd1669: RELPAGE <= 12'd555;
            12'd1670: RELPAGE <= 12'd1077;
            12'd1671: RELPAGE <= 12'd1599;
            12'd1672: RELPAGE <= 12'd68;
            12'd1673: RELPAGE <= 12'd590;
            12'd1674: RELPAGE <= 12'd1112;
            12'd1675: RELPAGE <= 12'd1634;
            12'd1676: RELPAGE <= 12'd103;
            12'd1677: RELPAGE <= 12'd625;
            12'd1678: RELPAGE <= 12'd1147;
            12'd1679: RELPAGE <= 12'd1669;
            12'd1680: RELPAGE <= 12'd138;
            12'd1681: RELPAGE <= 12'd660;
            12'd1682: RELPAGE <= 12'd1182;
            12'd1683: RELPAGE <= 12'd1704;
            12'd1684: RELPAGE <= 12'd173;
            12'd1685: RELPAGE <= 12'd695;
            12'd1686: RELPAGE <= 12'd1217;
            12'd1687: RELPAGE <= 12'd1739;
            12'd1688: RELPAGE <= 12'd208;
            12'd1689: RELPAGE <= 12'd730;
            12'd1690: RELPAGE <= 12'd1252;
            12'd1691: RELPAGE <= 12'd1774;
            12'd1692: RELPAGE <= 12'd243;
            12'd1693: RELPAGE <= 12'd765;
            12'd1694: RELPAGE <= 12'd1287;
            12'd1695: RELPAGE <= 12'd1809;
            12'd1696: RELPAGE <= 12'd278;
            12'd1697: RELPAGE <= 12'd800;
            12'd1698: RELPAGE <= 12'd1322;
            12'd1699: RELPAGE <= 12'd1844;
            12'd1700: RELPAGE <= 12'd313;
            12'd1701: RELPAGE <= 12'd835;
            12'd1702: RELPAGE <= 12'd1357;
            12'd1703: RELPAGE <= 12'd1879;
            12'd1704: RELPAGE <= 12'd348;
            12'd1705: RELPAGE <= 12'd870;
            12'd1706: RELPAGE <= 12'd1392;
            12'd1707: RELPAGE <= 12'd1914;
            12'd1708: RELPAGE <= 12'd383;
            12'd1709: RELPAGE <= 12'd905;
            12'd1710: RELPAGE <= 12'd1427;
            12'd1711: RELPAGE <= 12'd1949;
            12'd1712: RELPAGE <= 12'd418;
            12'd1713: RELPAGE <= 12'd940;
            12'd1714: RELPAGE <= 12'd1462;
            12'd1715: RELPAGE <= 12'd1984;
            12'd1716: RELPAGE <= 12'd453;
            12'd1717: RELPAGE <= 12'd975;
            12'd1718: RELPAGE <= 12'd1497;
            12'd1719: RELPAGE <= 12'd2019;
            12'd1720: RELPAGE <= 12'd488;
            12'd1721: RELPAGE <= 12'd1010;
            12'd1722: RELPAGE <= 12'd1532;
            12'd1723: RELPAGE <= 12'd1;
            12'd1724: RELPAGE <= 12'd523;
            12'd1725: RELPAGE <= 12'd1045;
            12'd1726: RELPAGE <= 12'd1567;
            12'd1727: RELPAGE <= 12'd36;
            12'd1728: RELPAGE <= 12'd558;
            12'd1729: RELPAGE <= 12'd1080;
            12'd1730: RELPAGE <= 12'd1602;
            12'd1731: RELPAGE <= 12'd71;
            12'd1732: RELPAGE <= 12'd593;
            12'd1733: RELPAGE <= 12'd1115;
            12'd1734: RELPAGE <= 12'd1637;
            12'd1735: RELPAGE <= 12'd106;
            12'd1736: RELPAGE <= 12'd628;
            12'd1737: RELPAGE <= 12'd1150;
            12'd1738: RELPAGE <= 12'd1672;
            12'd1739: RELPAGE <= 12'd141;
            12'd1740: RELPAGE <= 12'd663;
            12'd1741: RELPAGE <= 12'd1185;
            12'd1742: RELPAGE <= 12'd1707;
            12'd1743: RELPAGE <= 12'd176;
            12'd1744: RELPAGE <= 12'd698;
            12'd1745: RELPAGE <= 12'd1220;
            12'd1746: RELPAGE <= 12'd1742;
            12'd1747: RELPAGE <= 12'd211;
            12'd1748: RELPAGE <= 12'd733;
            12'd1749: RELPAGE <= 12'd1255;
            12'd1750: RELPAGE <= 12'd1777;
            12'd1751: RELPAGE <= 12'd246;
            12'd1752: RELPAGE <= 12'd768;
            12'd1753: RELPAGE <= 12'd1290;
            12'd1754: RELPAGE <= 12'd1812;
            12'd1755: RELPAGE <= 12'd281;
            12'd1756: RELPAGE <= 12'd803;
            12'd1757: RELPAGE <= 12'd1325;
            12'd1758: RELPAGE <= 12'd1847;
            12'd1759: RELPAGE <= 12'd316;
            12'd1760: RELPAGE <= 12'd838;
            12'd1761: RELPAGE <= 12'd1360;
            12'd1762: RELPAGE <= 12'd1882;
            12'd1763: RELPAGE <= 12'd351;
            12'd1764: RELPAGE <= 12'd873;
            12'd1765: RELPAGE <= 12'd1395;
            12'd1766: RELPAGE <= 12'd1917;
            12'd1767: RELPAGE <= 12'd386;
            12'd1768: RELPAGE <= 12'd908;
            12'd1769: RELPAGE <= 12'd1430;
            12'd1770: RELPAGE <= 12'd1952;
            12'd1771: RELPAGE <= 12'd421;
            12'd1772: RELPAGE <= 12'd943;
            12'd1773: RELPAGE <= 12'd1465;
            12'd1774: RELPAGE <= 12'd1987;
            12'd1775: RELPAGE <= 12'd456;
            12'd1776: RELPAGE <= 12'd978;
            12'd1777: RELPAGE <= 12'd1500;
            12'd1778: RELPAGE <= 12'd2022;
            12'd1779: RELPAGE <= 12'd491;
            12'd1780: RELPAGE <= 12'd1013;
            12'd1781: RELPAGE <= 12'd1535;
            12'd1782: RELPAGE <= 12'd4;
            12'd1783: RELPAGE <= 12'd526;
            12'd1784: RELPAGE <= 12'd1048;
            12'd1785: RELPAGE <= 12'd1570;
            12'd1786: RELPAGE <= 12'd39;
            12'd1787: RELPAGE <= 12'd561;
            12'd1788: RELPAGE <= 12'd1083;
            12'd1789: RELPAGE <= 12'd1605;
            12'd1790: RELPAGE <= 12'd74;
            12'd1791: RELPAGE <= 12'd596;
            12'd1792: RELPAGE <= 12'd1118;
            12'd1793: RELPAGE <= 12'd1640;
            12'd1794: RELPAGE <= 12'd109;
            12'd1795: RELPAGE <= 12'd631;
            12'd1796: RELPAGE <= 12'd1153;
            12'd1797: RELPAGE <= 12'd1675;
            12'd1798: RELPAGE <= 12'd144;
            12'd1799: RELPAGE <= 12'd666;
            12'd1800: RELPAGE <= 12'd1188;
            12'd1801: RELPAGE <= 12'd1710;
            12'd1802: RELPAGE <= 12'd179;
            12'd1803: RELPAGE <= 12'd701;
            12'd1804: RELPAGE <= 12'd1223;
            12'd1805: RELPAGE <= 12'd1745;
            12'd1806: RELPAGE <= 12'd214;
            12'd1807: RELPAGE <= 12'd736;
            12'd1808: RELPAGE <= 12'd1258;
            12'd1809: RELPAGE <= 12'd1780;
            12'd1810: RELPAGE <= 12'd249;
            12'd1811: RELPAGE <= 12'd771;
            12'd1812: RELPAGE <= 12'd1293;
            12'd1813: RELPAGE <= 12'd1815;
            12'd1814: RELPAGE <= 12'd284;
            12'd1815: RELPAGE <= 12'd806;
            12'd1816: RELPAGE <= 12'd1328;
            12'd1817: RELPAGE <= 12'd1850;
            12'd1818: RELPAGE <= 12'd319;
            12'd1819: RELPAGE <= 12'd841;
            12'd1820: RELPAGE <= 12'd1363;
            12'd1821: RELPAGE <= 12'd1885;
            12'd1822: RELPAGE <= 12'd354;
            12'd1823: RELPAGE <= 12'd876;
            12'd1824: RELPAGE <= 12'd1398;
            12'd1825: RELPAGE <= 12'd1920;
            12'd1826: RELPAGE <= 12'd389;
            12'd1827: RELPAGE <= 12'd911;
            12'd1828: RELPAGE <= 12'd1433;
            12'd1829: RELPAGE <= 12'd1955;
            12'd1830: RELPAGE <= 12'd424;
            12'd1831: RELPAGE <= 12'd946;
            12'd1832: RELPAGE <= 12'd1468;
            12'd1833: RELPAGE <= 12'd1990;
            12'd1834: RELPAGE <= 12'd459;
            12'd1835: RELPAGE <= 12'd981;
            12'd1836: RELPAGE <= 12'd1503;
            12'd1837: RELPAGE <= 12'd2025;
            12'd1838: RELPAGE <= 12'd494;
            12'd1839: RELPAGE <= 12'd1016;
            12'd1840: RELPAGE <= 12'd1538;
            12'd1841: RELPAGE <= 12'd7;
            12'd1842: RELPAGE <= 12'd529;
            12'd1843: RELPAGE <= 12'd1051;
            12'd1844: RELPAGE <= 12'd1573;
            12'd1845: RELPAGE <= 12'd42;
            12'd1846: RELPAGE <= 12'd564;
            12'd1847: RELPAGE <= 12'd1086;
            12'd1848: RELPAGE <= 12'd1608;
            12'd1849: RELPAGE <= 12'd77;
            12'd1850: RELPAGE <= 12'd599;
            12'd1851: RELPAGE <= 12'd1121;
            12'd1852: RELPAGE <= 12'd1643;
            12'd1853: RELPAGE <= 12'd112;
            12'd1854: RELPAGE <= 12'd634;
            12'd1855: RELPAGE <= 12'd1156;
            12'd1856: RELPAGE <= 12'd1678;
            12'd1857: RELPAGE <= 12'd147;
            12'd1858: RELPAGE <= 12'd669;
            12'd1859: RELPAGE <= 12'd1191;
            12'd1860: RELPAGE <= 12'd1713;
            12'd1861: RELPAGE <= 12'd182;
            12'd1862: RELPAGE <= 12'd704;
            12'd1863: RELPAGE <= 12'd1226;
            12'd1864: RELPAGE <= 12'd1748;
            12'd1865: RELPAGE <= 12'd217;
            12'd1866: RELPAGE <= 12'd739;
            12'd1867: RELPAGE <= 12'd1261;
            12'd1868: RELPAGE <= 12'd1783;
            12'd1869: RELPAGE <= 12'd252;
            12'd1870: RELPAGE <= 12'd774;
            12'd1871: RELPAGE <= 12'd1296;
            12'd1872: RELPAGE <= 12'd1818;
            12'd1873: RELPAGE <= 12'd287;
            12'd1874: RELPAGE <= 12'd809;
            12'd1875: RELPAGE <= 12'd1331;
            12'd1876: RELPAGE <= 12'd1853;
            12'd1877: RELPAGE <= 12'd322;
            12'd1878: RELPAGE <= 12'd844;
            12'd1879: RELPAGE <= 12'd1366;
            12'd1880: RELPAGE <= 12'd1888;
            12'd1881: RELPAGE <= 12'd357;
            12'd1882: RELPAGE <= 12'd879;
            12'd1883: RELPAGE <= 12'd1401;
            12'd1884: RELPAGE <= 12'd1923;
            12'd1885: RELPAGE <= 12'd392;
            12'd1886: RELPAGE <= 12'd914;
            12'd1887: RELPAGE <= 12'd1436;
            12'd1888: RELPAGE <= 12'd1958;
            12'd1889: RELPAGE <= 12'd427;
            12'd1890: RELPAGE <= 12'd949;
            12'd1891: RELPAGE <= 12'd1471;
            12'd1892: RELPAGE <= 12'd1993;
            12'd1893: RELPAGE <= 12'd462;
            12'd1894: RELPAGE <= 12'd984;
            12'd1895: RELPAGE <= 12'd1506;
            12'd1896: RELPAGE <= 12'd2028;
            12'd1897: RELPAGE <= 12'd497;
            12'd1898: RELPAGE <= 12'd1019;
            12'd1899: RELPAGE <= 12'd1541;
            12'd1900: RELPAGE <= 12'd10;
            12'd1901: RELPAGE <= 12'd532;
            12'd1902: RELPAGE <= 12'd1054;
            12'd1903: RELPAGE <= 12'd1576;
            12'd1904: RELPAGE <= 12'd45;
            12'd1905: RELPAGE <= 12'd567;
            12'd1906: RELPAGE <= 12'd1089;
            12'd1907: RELPAGE <= 12'd1611;
            12'd1908: RELPAGE <= 12'd80;
            12'd1909: RELPAGE <= 12'd602;
            12'd1910: RELPAGE <= 12'd1124;
            12'd1911: RELPAGE <= 12'd1646;
            12'd1912: RELPAGE <= 12'd115;
            12'd1913: RELPAGE <= 12'd637;
            12'd1914: RELPAGE <= 12'd1159;
            12'd1915: RELPAGE <= 12'd1681;
            12'd1916: RELPAGE <= 12'd150;
            12'd1917: RELPAGE <= 12'd672;
            12'd1918: RELPAGE <= 12'd1194;
            12'd1919: RELPAGE <= 12'd1716;
            12'd1920: RELPAGE <= 12'd185;
            12'd1921: RELPAGE <= 12'd707;
            12'd1922: RELPAGE <= 12'd1229;
            12'd1923: RELPAGE <= 12'd1751;
            12'd1924: RELPAGE <= 12'd220;
            12'd1925: RELPAGE <= 12'd742;
            12'd1926: RELPAGE <= 12'd1264;
            12'd1927: RELPAGE <= 12'd1786;
            12'd1928: RELPAGE <= 12'd255;
            12'd1929: RELPAGE <= 12'd777;
            12'd1930: RELPAGE <= 12'd1299;
            12'd1931: RELPAGE <= 12'd1821;
            12'd1932: RELPAGE <= 12'd290;
            12'd1933: RELPAGE <= 12'd812;
            12'd1934: RELPAGE <= 12'd1334;
            12'd1935: RELPAGE <= 12'd1856;
            12'd1936: RELPAGE <= 12'd325;
            12'd1937: RELPAGE <= 12'd847;
            12'd1938: RELPAGE <= 12'd1369;
            12'd1939: RELPAGE <= 12'd1891;
            12'd1940: RELPAGE <= 12'd360;
            12'd1941: RELPAGE <= 12'd882;
            12'd1942: RELPAGE <= 12'd1404;
            12'd1943: RELPAGE <= 12'd1926;
            12'd1944: RELPAGE <= 12'd395;
            12'd1945: RELPAGE <= 12'd917;
            12'd1946: RELPAGE <= 12'd1439;
            12'd1947: RELPAGE <= 12'd1961;
            12'd1948: RELPAGE <= 12'd430;
            12'd1949: RELPAGE <= 12'd952;
            12'd1950: RELPAGE <= 12'd1474;
            12'd1951: RELPAGE <= 12'd1996;
            12'd1952: RELPAGE <= 12'd465;
            12'd1953: RELPAGE <= 12'd987;
            12'd1954: RELPAGE <= 12'd1509;
            12'd1955: RELPAGE <= 12'd2031;
            12'd1956: RELPAGE <= 12'd500;
            12'd1957: RELPAGE <= 12'd1022;
            12'd1958: RELPAGE <= 12'd1544;
            12'd1959: RELPAGE <= 12'd13;
            12'd1960: RELPAGE <= 12'd535;
            12'd1961: RELPAGE <= 12'd1057;
            12'd1962: RELPAGE <= 12'd1579;
            12'd1963: RELPAGE <= 12'd48;
            12'd1964: RELPAGE <= 12'd570;
            12'd1965: RELPAGE <= 12'd1092;
            12'd1966: RELPAGE <= 12'd1614;
            12'd1967: RELPAGE <= 12'd83;
            12'd1968: RELPAGE <= 12'd605;
            12'd1969: RELPAGE <= 12'd1127;
            12'd1970: RELPAGE <= 12'd1649;
            12'd1971: RELPAGE <= 12'd118;
            12'd1972: RELPAGE <= 12'd640;
            12'd1973: RELPAGE <= 12'd1162;
            12'd1974: RELPAGE <= 12'd1684;
            12'd1975: RELPAGE <= 12'd153;
            12'd1976: RELPAGE <= 12'd675;
            12'd1977: RELPAGE <= 12'd1197;
            12'd1978: RELPAGE <= 12'd1719;
            12'd1979: RELPAGE <= 12'd188;
            12'd1980: RELPAGE <= 12'd710;
            12'd1981: RELPAGE <= 12'd1232;
            12'd1982: RELPAGE <= 12'd1754;
            12'd1983: RELPAGE <= 12'd223;
            12'd1984: RELPAGE <= 12'd745;
            12'd1985: RELPAGE <= 12'd1267;
            12'd1986: RELPAGE <= 12'd1789;
            12'd1987: RELPAGE <= 12'd258;
            12'd1988: RELPAGE <= 12'd780;
            12'd1989: RELPAGE <= 12'd1302;
            12'd1990: RELPAGE <= 12'd1824;
            12'd1991: RELPAGE <= 12'd293;
            12'd1992: RELPAGE <= 12'd815;
            12'd1993: RELPAGE <= 12'd1337;
            12'd1994: RELPAGE <= 12'd1859;
            12'd1995: RELPAGE <= 12'd328;
            12'd1996: RELPAGE <= 12'd850;
            12'd1997: RELPAGE <= 12'd1372;
            12'd1998: RELPAGE <= 12'd1894;
            12'd1999: RELPAGE <= 12'd363;
            12'd2000: RELPAGE <= 12'd885;
            12'd2001: RELPAGE <= 12'd1407;
            12'd2002: RELPAGE <= 12'd1929;
            12'd2003: RELPAGE <= 12'd398;
            12'd2004: RELPAGE <= 12'd920;
            12'd2005: RELPAGE <= 12'd1442;
            12'd2006: RELPAGE <= 12'd1964;
            12'd2007: RELPAGE <= 12'd433;
            12'd2008: RELPAGE <= 12'd955;
            12'd2009: RELPAGE <= 12'd1477;
            12'd2010: RELPAGE <= 12'd1999;
            12'd2011: RELPAGE <= 12'd468;
            12'd2012: RELPAGE <= 12'd990;
            12'd2013: RELPAGE <= 12'd1512;
            12'd2014: RELPAGE <= 12'd2034;
            12'd2015: RELPAGE <= 12'd503;
            12'd2016: RELPAGE <= 12'd1025;
            12'd2017: RELPAGE <= 12'd1547;
            12'd2018: RELPAGE <= 12'd16;
            12'd2019: RELPAGE <= 12'd538;
            12'd2020: RELPAGE <= 12'd1060;
            12'd2021: RELPAGE <= 12'd1582;
            12'd2022: RELPAGE <= 12'd51;
            12'd2023: RELPAGE <= 12'd573;
            12'd2024: RELPAGE <= 12'd1095;
            12'd2025: RELPAGE <= 12'd1617;
            12'd2026: RELPAGE <= 12'd86;
            12'd2027: RELPAGE <= 12'd608;
            12'd2028: RELPAGE <= 12'd1130;
            12'd2029: RELPAGE <= 12'd1652;
            12'd2030: RELPAGE <= 12'd121;
            12'd2031: RELPAGE <= 12'd643;
            12'd2032: RELPAGE <= 12'd1165;
            12'd2033: RELPAGE <= 12'd1687;
            12'd2034: RELPAGE <= 12'd156;
            12'd2035: RELPAGE <= 12'd678;
            12'd2036: RELPAGE <= 12'd1200;
            12'd2037: RELPAGE <= 12'd1722;
            12'd2038: RELPAGE <= 12'd191;
            12'd2039: RELPAGE <= 12'd713;
            12'd2040: RELPAGE <= 12'd1235;
            12'd2041: RELPAGE <= 12'd1757;
            12'd2042: RELPAGE <= 12'd226;
            12'd2043: RELPAGE <= 12'd748;
            12'd2044: RELPAGE <= 12'd1270;
            12'd2045: RELPAGE <= 12'd1792;
            12'd2046: RELPAGE <= 12'd261;
            12'd2047: RELPAGE <= 12'd783;
            12'd2048: RELPAGE <= 12'd1305;
            12'd2049: RELPAGE <= 12'd1827;
            12'd2050: RELPAGE <= 12'd296;
            12'd2051: RELPAGE <= 12'd818;
            12'd2052: RELPAGE <= 12'd1340;
            12'd2053: RELPAGE <= 12'd1862;
            12'd2054: RELPAGE <= 12'd4095;
            12'd2055: RELPAGE <= 12'd4095;
            12'd2056: RELPAGE <= 12'd4095;
            12'd2057: RELPAGE <= 12'd4095;
            12'd2058: RELPAGE <= 12'd4095;
            12'd2059: RELPAGE <= 12'd4095;
            12'd2060: RELPAGE <= 12'd4095;
            12'd2061: RELPAGE <= 12'd4095;
            12'd2062: RELPAGE <= 12'd4095;
            12'd2063: RELPAGE <= 12'd4095;
            12'd2064: RELPAGE <= 12'd4095;
            12'd2065: RELPAGE <= 12'd4095;
            12'd2066: RELPAGE <= 12'd4095;
            12'd2067: RELPAGE <= 12'd4095;
            12'd2068: RELPAGE <= 12'd4095;
            12'd2069: RELPAGE <= 12'd4095;
            12'd2070: RELPAGE <= 12'd4095;
            12'd2071: RELPAGE <= 12'd4095;
            12'd2072: RELPAGE <= 12'd4095;
            12'd2073: RELPAGE <= 12'd4095;
            12'd2074: RELPAGE <= 12'd4095;
            12'd2075: RELPAGE <= 12'd4095;
            12'd2076: RELPAGE <= 12'd4095;
            12'd2077: RELPAGE <= 12'd4095;
            12'd2078: RELPAGE <= 12'd4095;
            12'd2079: RELPAGE <= 12'd4095;
            12'd2080: RELPAGE <= 12'd4095;
            12'd2081: RELPAGE <= 12'd4095;
            12'd2082: RELPAGE <= 12'd4095;
            12'd2083: RELPAGE <= 12'd4095;
            12'd2084: RELPAGE <= 12'd4095;
            12'd2085: RELPAGE <= 12'd4095;
            12'd2086: RELPAGE <= 12'd4095;
            12'd2087: RELPAGE <= 12'd4095;
            12'd2088: RELPAGE <= 12'd4095;
            12'd2089: RELPAGE <= 12'd4095;
            12'd2090: RELPAGE <= 12'd4095;
            12'd2091: RELPAGE <= 12'd4095;
            12'd2092: RELPAGE <= 12'd4095;
            12'd2093: RELPAGE <= 12'd4095;
            12'd2094: RELPAGE <= 12'd4095;
            12'd2095: RELPAGE <= 12'd4095;
            12'd2096: RELPAGE <= 12'd4095;
            12'd2097: RELPAGE <= 12'd4095;
            12'd2098: RELPAGE <= 12'd4095;
            12'd2099: RELPAGE <= 12'd4095;
            12'd2100: RELPAGE <= 12'd4095;
            12'd2101: RELPAGE <= 12'd4095;
            12'd2102: RELPAGE <= 12'd4095;
            12'd2103: RELPAGE <= 12'd4095;
            12'd2104: RELPAGE <= 12'd4095;
            12'd2105: RELPAGE <= 12'd4095;
            12'd2106: RELPAGE <= 12'd4095;
            12'd2107: RELPAGE <= 12'd4095;
            12'd2108: RELPAGE <= 12'd4095;
            12'd2109: RELPAGE <= 12'd4095;
            12'd2110: RELPAGE <= 12'd4095;
            12'd2111: RELPAGE <= 12'd4095;
            12'd2112: RELPAGE <= 12'd4095;
            12'd2113: RELPAGE <= 12'd4095;
            12'd2114: RELPAGE <= 12'd4095;
            12'd2115: RELPAGE <= 12'd4095;
            12'd2116: RELPAGE <= 12'd4095;
            12'd2117: RELPAGE <= 12'd4095;
            12'd2118: RELPAGE <= 12'd4095;
            12'd2119: RELPAGE <= 12'd4095;
            12'd2120: RELPAGE <= 12'd4095;
            12'd2121: RELPAGE <= 12'd4095;
            12'd2122: RELPAGE <= 12'd4095;
            12'd2123: RELPAGE <= 12'd4095;
            12'd2124: RELPAGE <= 12'd4095;
            12'd2125: RELPAGE <= 12'd4095;
            12'd2126: RELPAGE <= 12'd4095;
            12'd2127: RELPAGE <= 12'd4095;
            12'd2128: RELPAGE <= 12'd4095;
            12'd2129: RELPAGE <= 12'd4095;
            12'd2130: RELPAGE <= 12'd4095;
            12'd2131: RELPAGE <= 12'd4095;
            12'd2132: RELPAGE <= 12'd4095;
            12'd2133: RELPAGE <= 12'd4095;
            12'd2134: RELPAGE <= 12'd4095;
            12'd2135: RELPAGE <= 12'd4095;
            12'd2136: RELPAGE <= 12'd4095;
            12'd2137: RELPAGE <= 12'd4095;
            12'd2138: RELPAGE <= 12'd4095;
            12'd2139: RELPAGE <= 12'd4095;
            12'd2140: RELPAGE <= 12'd4095;
            12'd2141: RELPAGE <= 12'd4095;
            12'd2142: RELPAGE <= 12'd4095;
            12'd2143: RELPAGE <= 12'd4095;
            12'd2144: RELPAGE <= 12'd4095;
            12'd2145: RELPAGE <= 12'd4095;
            12'd2146: RELPAGE <= 12'd4095;
            12'd2147: RELPAGE <= 12'd4095;
            12'd2148: RELPAGE <= 12'd4095;
            12'd2149: RELPAGE <= 12'd4095;
            12'd2150: RELPAGE <= 12'd4095;
            12'd2151: RELPAGE <= 12'd4095;
            12'd2152: RELPAGE <= 12'd4095;
            12'd2153: RELPAGE <= 12'd4095;
            12'd2154: RELPAGE <= 12'd4095;
            12'd2155: RELPAGE <= 12'd4095;
            12'd2156: RELPAGE <= 12'd4095;
            12'd2157: RELPAGE <= 12'd4095;
            12'd2158: RELPAGE <= 12'd4095;
            12'd2159: RELPAGE <= 12'd4095;
            12'd2160: RELPAGE <= 12'd4095;
            12'd2161: RELPAGE <= 12'd4095;
            12'd2162: RELPAGE <= 12'd4095;
            12'd2163: RELPAGE <= 12'd4095;
            12'd2164: RELPAGE <= 12'd4095;
            12'd2165: RELPAGE <= 12'd4095;
            12'd2166: RELPAGE <= 12'd4095;
            12'd2167: RELPAGE <= 12'd4095;
            12'd2168: RELPAGE <= 12'd4095;
            12'd2169: RELPAGE <= 12'd4095;
            12'd2170: RELPAGE <= 12'd4095;
            12'd2171: RELPAGE <= 12'd4095;
            12'd2172: RELPAGE <= 12'd4095;
            12'd2173: RELPAGE <= 12'd4095;
            12'd2174: RELPAGE <= 12'd4095;
            12'd2175: RELPAGE <= 12'd4095;
            12'd2176: RELPAGE <= 12'd4095;
            12'd2177: RELPAGE <= 12'd4095;
            12'd2178: RELPAGE <= 12'd4095;
            12'd2179: RELPAGE <= 12'd4095;
            12'd2180: RELPAGE <= 12'd4095;
            12'd2181: RELPAGE <= 12'd4095;
            12'd2182: RELPAGE <= 12'd4095;
            12'd2183: RELPAGE <= 12'd4095;
            12'd2184: RELPAGE <= 12'd4095;
            12'd2185: RELPAGE <= 12'd4095;
            12'd2186: RELPAGE <= 12'd4095;
            12'd2187: RELPAGE <= 12'd4095;
            12'd2188: RELPAGE <= 12'd4095;
            12'd2189: RELPAGE <= 12'd4095;
            12'd2190: RELPAGE <= 12'd4095;
            12'd2191: RELPAGE <= 12'd4095;
            12'd2192: RELPAGE <= 12'd4095;
            12'd2193: RELPAGE <= 12'd4095;
            12'd2194: RELPAGE <= 12'd4095;
            12'd2195: RELPAGE <= 12'd4095;
            12'd2196: RELPAGE <= 12'd4095;
            12'd2197: RELPAGE <= 12'd4095;
            12'd2198: RELPAGE <= 12'd4095;
            12'd2199: RELPAGE <= 12'd4095;
            12'd2200: RELPAGE <= 12'd4095;
            12'd2201: RELPAGE <= 12'd4095;
            12'd2202: RELPAGE <= 12'd4095;
            12'd2203: RELPAGE <= 12'd4095;
            12'd2204: RELPAGE <= 12'd4095;
            12'd2205: RELPAGE <= 12'd4095;
            12'd2206: RELPAGE <= 12'd4095;
            12'd2207: RELPAGE <= 12'd4095;
            12'd2208: RELPAGE <= 12'd4095;
            12'd2209: RELPAGE <= 12'd4095;
            12'd2210: RELPAGE <= 12'd4095;
            12'd2211: RELPAGE <= 12'd4095;
            12'd2212: RELPAGE <= 12'd4095;
            12'd2213: RELPAGE <= 12'd4095;
            12'd2214: RELPAGE <= 12'd4095;
            12'd2215: RELPAGE <= 12'd4095;
            12'd2216: RELPAGE <= 12'd4095;
            12'd2217: RELPAGE <= 12'd4095;
            12'd2218: RELPAGE <= 12'd4095;
            12'd2219: RELPAGE <= 12'd4095;
            12'd2220: RELPAGE <= 12'd4095;
            12'd2221: RELPAGE <= 12'd4095;
            12'd2222: RELPAGE <= 12'd4095;
            12'd2223: RELPAGE <= 12'd4095;
            12'd2224: RELPAGE <= 12'd4095;
            12'd2225: RELPAGE <= 12'd4095;
            12'd2226: RELPAGE <= 12'd4095;
            12'd2227: RELPAGE <= 12'd4095;
            12'd2228: RELPAGE <= 12'd4095;
            12'd2229: RELPAGE <= 12'd4095;
            12'd2230: RELPAGE <= 12'd4095;
            12'd2231: RELPAGE <= 12'd4095;
            12'd2232: RELPAGE <= 12'd4095;
            12'd2233: RELPAGE <= 12'd4095;
            12'd2234: RELPAGE <= 12'd4095;
            12'd2235: RELPAGE <= 12'd4095;
            12'd2236: RELPAGE <= 12'd4095;
            12'd2237: RELPAGE <= 12'd4095;
            12'd2238: RELPAGE <= 12'd4095;
            12'd2239: RELPAGE <= 12'd4095;
            12'd2240: RELPAGE <= 12'd4095;
            12'd2241: RELPAGE <= 12'd4095;
            12'd2242: RELPAGE <= 12'd4095;
            12'd2243: RELPAGE <= 12'd4095;
            12'd2244: RELPAGE <= 12'd4095;
            12'd2245: RELPAGE <= 12'd4095;
            12'd2246: RELPAGE <= 12'd4095;
            12'd2247: RELPAGE <= 12'd4095;
            12'd2248: RELPAGE <= 12'd4095;
            12'd2249: RELPAGE <= 12'd4095;
            12'd2250: RELPAGE <= 12'd4095;
            12'd2251: RELPAGE <= 12'd4095;
            12'd2252: RELPAGE <= 12'd4095;
            12'd2253: RELPAGE <= 12'd4095;
            12'd2254: RELPAGE <= 12'd4095;
            12'd2255: RELPAGE <= 12'd4095;
            12'd2256: RELPAGE <= 12'd4095;
            12'd2257: RELPAGE <= 12'd4095;
            12'd2258: RELPAGE <= 12'd4095;
            12'd2259: RELPAGE <= 12'd4095;
            12'd2260: RELPAGE <= 12'd4095;
            12'd2261: RELPAGE <= 12'd4095;
            12'd2262: RELPAGE <= 12'd4095;
            12'd2263: RELPAGE <= 12'd4095;
            12'd2264: RELPAGE <= 12'd4095;
            12'd2265: RELPAGE <= 12'd4095;
            12'd2266: RELPAGE <= 12'd4095;
            12'd2267: RELPAGE <= 12'd4095;
            12'd2268: RELPAGE <= 12'd4095;
            12'd2269: RELPAGE <= 12'd4095;
            12'd2270: RELPAGE <= 12'd4095;
            12'd2271: RELPAGE <= 12'd4095;
            12'd2272: RELPAGE <= 12'd4095;
            12'd2273: RELPAGE <= 12'd4095;
            12'd2274: RELPAGE <= 12'd4095;
            12'd2275: RELPAGE <= 12'd4095;
            12'd2276: RELPAGE <= 12'd4095;
            12'd2277: RELPAGE <= 12'd4095;
            12'd2278: RELPAGE <= 12'd4095;
            12'd2279: RELPAGE <= 12'd4095;
            12'd2280: RELPAGE <= 12'd4095;
            12'd2281: RELPAGE <= 12'd4095;
            12'd2282: RELPAGE <= 12'd4095;
            12'd2283: RELPAGE <= 12'd4095;
            12'd2284: RELPAGE <= 12'd4095;
            12'd2285: RELPAGE <= 12'd4095;
            12'd2286: RELPAGE <= 12'd4095;
            12'd2287: RELPAGE <= 12'd4095;
            12'd2288: RELPAGE <= 12'd4095;
            12'd2289: RELPAGE <= 12'd4095;
            12'd2290: RELPAGE <= 12'd4095;
            12'd2291: RELPAGE <= 12'd4095;
            12'd2292: RELPAGE <= 12'd4095;
            12'd2293: RELPAGE <= 12'd4095;
            12'd2294: RELPAGE <= 12'd4095;
            12'd2295: RELPAGE <= 12'd4095;
            12'd2296: RELPAGE <= 12'd4095;
            12'd2297: RELPAGE <= 12'd4095;
            12'd2298: RELPAGE <= 12'd4095;
            12'd2299: RELPAGE <= 12'd4095;
            12'd2300: RELPAGE <= 12'd4095;
            12'd2301: RELPAGE <= 12'd4095;
            12'd2302: RELPAGE <= 12'd4095;
            12'd2303: RELPAGE <= 12'd4095;
            12'd2304: RELPAGE <= 12'd4095;
            12'd2305: RELPAGE <= 12'd4095;
            12'd2306: RELPAGE <= 12'd4095;
            12'd2307: RELPAGE <= 12'd4095;
            12'd2308: RELPAGE <= 12'd4095;
            12'd2309: RELPAGE <= 12'd4095;
            12'd2310: RELPAGE <= 12'd4095;
            12'd2311: RELPAGE <= 12'd4095;
            12'd2312: RELPAGE <= 12'd4095;
            12'd2313: RELPAGE <= 12'd4095;
            12'd2314: RELPAGE <= 12'd4095;
            12'd2315: RELPAGE <= 12'd4095;
            12'd2316: RELPAGE <= 12'd4095;
            12'd2317: RELPAGE <= 12'd4095;
            12'd2318: RELPAGE <= 12'd4095;
            12'd2319: RELPAGE <= 12'd4095;
            12'd2320: RELPAGE <= 12'd4095;
            12'd2321: RELPAGE <= 12'd4095;
            12'd2322: RELPAGE <= 12'd4095;
            12'd2323: RELPAGE <= 12'd4095;
            12'd2324: RELPAGE <= 12'd4095;
            12'd2325: RELPAGE <= 12'd4095;
            12'd2326: RELPAGE <= 12'd4095;
            12'd2327: RELPAGE <= 12'd4095;
            12'd2328: RELPAGE <= 12'd4095;
            12'd2329: RELPAGE <= 12'd4095;
            12'd2330: RELPAGE <= 12'd4095;
            12'd2331: RELPAGE <= 12'd4095;
            12'd2332: RELPAGE <= 12'd4095;
            12'd2333: RELPAGE <= 12'd4095;
            12'd2334: RELPAGE <= 12'd4095;
            12'd2335: RELPAGE <= 12'd4095;
            12'd2336: RELPAGE <= 12'd4095;
            12'd2337: RELPAGE <= 12'd4095;
            12'd2338: RELPAGE <= 12'd4095;
            12'd2339: RELPAGE <= 12'd4095;
            12'd2340: RELPAGE <= 12'd4095;
            12'd2341: RELPAGE <= 12'd4095;
            12'd2342: RELPAGE <= 12'd4095;
            12'd2343: RELPAGE <= 12'd4095;
            12'd2344: RELPAGE <= 12'd4095;
            12'd2345: RELPAGE <= 12'd4095;
            12'd2346: RELPAGE <= 12'd4095;
            12'd2347: RELPAGE <= 12'd4095;
            12'd2348: RELPAGE <= 12'd4095;
            12'd2349: RELPAGE <= 12'd4095;
            12'd2350: RELPAGE <= 12'd4095;
            12'd2351: RELPAGE <= 12'd4095;
            12'd2352: RELPAGE <= 12'd4095;
            12'd2353: RELPAGE <= 12'd4095;
            12'd2354: RELPAGE <= 12'd4095;
            12'd2355: RELPAGE <= 12'd4095;
            12'd2356: RELPAGE <= 12'd4095;
            12'd2357: RELPAGE <= 12'd4095;
            12'd2358: RELPAGE <= 12'd4095;
            12'd2359: RELPAGE <= 12'd4095;
            12'd2360: RELPAGE <= 12'd4095;
            12'd2361: RELPAGE <= 12'd4095;
            12'd2362: RELPAGE <= 12'd4095;
            12'd2363: RELPAGE <= 12'd4095;
            12'd2364: RELPAGE <= 12'd4095;
            12'd2365: RELPAGE <= 12'd4095;
            12'd2366: RELPAGE <= 12'd4095;
            12'd2367: RELPAGE <= 12'd4095;
            12'd2368: RELPAGE <= 12'd4095;
            12'd2369: RELPAGE <= 12'd4095;
            12'd2370: RELPAGE <= 12'd4095;
            12'd2371: RELPAGE <= 12'd4095;
            12'd2372: RELPAGE <= 12'd4095;
            12'd2373: RELPAGE <= 12'd4095;
            12'd2374: RELPAGE <= 12'd4095;
            12'd2375: RELPAGE <= 12'd4095;
            12'd2376: RELPAGE <= 12'd4095;
            12'd2377: RELPAGE <= 12'd4095;
            12'd2378: RELPAGE <= 12'd4095;
            12'd2379: RELPAGE <= 12'd4095;
            12'd2380: RELPAGE <= 12'd4095;
            12'd2381: RELPAGE <= 12'd4095;
            12'd2382: RELPAGE <= 12'd4095;
            12'd2383: RELPAGE <= 12'd4095;
            12'd2384: RELPAGE <= 12'd4095;
            12'd2385: RELPAGE <= 12'd4095;
            12'd2386: RELPAGE <= 12'd4095;
            12'd2387: RELPAGE <= 12'd4095;
            12'd2388: RELPAGE <= 12'd4095;
            12'd2389: RELPAGE <= 12'd4095;
            12'd2390: RELPAGE <= 12'd4095;
            12'd2391: RELPAGE <= 12'd4095;
            12'd2392: RELPAGE <= 12'd4095;
            12'd2393: RELPAGE <= 12'd4095;
            12'd2394: RELPAGE <= 12'd4095;
            12'd2395: RELPAGE <= 12'd4095;
            12'd2396: RELPAGE <= 12'd4095;
            12'd2397: RELPAGE <= 12'd4095;
            12'd2398: RELPAGE <= 12'd4095;
            12'd2399: RELPAGE <= 12'd4095;
            12'd2400: RELPAGE <= 12'd4095;
            12'd2401: RELPAGE <= 12'd4095;
            12'd2402: RELPAGE <= 12'd4095;
            12'd2403: RELPAGE <= 12'd4095;
            12'd2404: RELPAGE <= 12'd4095;
            12'd2405: RELPAGE <= 12'd4095;
            12'd2406: RELPAGE <= 12'd4095;
            12'd2407: RELPAGE <= 12'd4095;
            12'd2408: RELPAGE <= 12'd4095;
            12'd2409: RELPAGE <= 12'd4095;
            12'd2410: RELPAGE <= 12'd4095;
            12'd2411: RELPAGE <= 12'd4095;
            12'd2412: RELPAGE <= 12'd4095;
            12'd2413: RELPAGE <= 12'd4095;
            12'd2414: RELPAGE <= 12'd4095;
            12'd2415: RELPAGE <= 12'd4095;
            12'd2416: RELPAGE <= 12'd4095;
            12'd2417: RELPAGE <= 12'd4095;
            12'd2418: RELPAGE <= 12'd4095;
            12'd2419: RELPAGE <= 12'd4095;
            12'd2420: RELPAGE <= 12'd4095;
            12'd2421: RELPAGE <= 12'd4095;
            12'd2422: RELPAGE <= 12'd4095;
            12'd2423: RELPAGE <= 12'd4095;
            12'd2424: RELPAGE <= 12'd4095;
            12'd2425: RELPAGE <= 12'd4095;
            12'd2426: RELPAGE <= 12'd4095;
            12'd2427: RELPAGE <= 12'd4095;
            12'd2428: RELPAGE <= 12'd4095;
            12'd2429: RELPAGE <= 12'd4095;
            12'd2430: RELPAGE <= 12'd4095;
            12'd2431: RELPAGE <= 12'd4095;
            12'd2432: RELPAGE <= 12'd4095;
            12'd2433: RELPAGE <= 12'd4095;
            12'd2434: RELPAGE <= 12'd4095;
            12'd2435: RELPAGE <= 12'd4095;
            12'd2436: RELPAGE <= 12'd4095;
            12'd2437: RELPAGE <= 12'd4095;
            12'd2438: RELPAGE <= 12'd4095;
            12'd2439: RELPAGE <= 12'd4095;
            12'd2440: RELPAGE <= 12'd4095;
            12'd2441: RELPAGE <= 12'd4095;
            12'd2442: RELPAGE <= 12'd4095;
            12'd2443: RELPAGE <= 12'd4095;
            12'd2444: RELPAGE <= 12'd4095;
            12'd2445: RELPAGE <= 12'd4095;
            12'd2446: RELPAGE <= 12'd4095;
            12'd2447: RELPAGE <= 12'd4095;
            12'd2448: RELPAGE <= 12'd4095;
            12'd2449: RELPAGE <= 12'd4095;
            12'd2450: RELPAGE <= 12'd4095;
            12'd2451: RELPAGE <= 12'd4095;
            12'd2452: RELPAGE <= 12'd4095;
            12'd2453: RELPAGE <= 12'd4095;
            12'd2454: RELPAGE <= 12'd4095;
            12'd2455: RELPAGE <= 12'd4095;
            12'd2456: RELPAGE <= 12'd4095;
            12'd2457: RELPAGE <= 12'd4095;
            12'd2458: RELPAGE <= 12'd4095;
            12'd2459: RELPAGE <= 12'd4095;
            12'd2460: RELPAGE <= 12'd4095;
            12'd2461: RELPAGE <= 12'd4095;
            12'd2462: RELPAGE <= 12'd4095;
            12'd2463: RELPAGE <= 12'd4095;
            12'd2464: RELPAGE <= 12'd4095;
            12'd2465: RELPAGE <= 12'd4095;
            12'd2466: RELPAGE <= 12'd4095;
            12'd2467: RELPAGE <= 12'd4095;
            12'd2468: RELPAGE <= 12'd4095;
            12'd2469: RELPAGE <= 12'd4095;
            12'd2470: RELPAGE <= 12'd4095;
            12'd2471: RELPAGE <= 12'd4095;
            12'd2472: RELPAGE <= 12'd4095;
            12'd2473: RELPAGE <= 12'd4095;
            12'd2474: RELPAGE <= 12'd4095;
            12'd2475: RELPAGE <= 12'd4095;
            12'd2476: RELPAGE <= 12'd4095;
            12'd2477: RELPAGE <= 12'd4095;
            12'd2478: RELPAGE <= 12'd4095;
            12'd2479: RELPAGE <= 12'd4095;
            12'd2480: RELPAGE <= 12'd4095;
            12'd2481: RELPAGE <= 12'd4095;
            12'd2482: RELPAGE <= 12'd4095;
            12'd2483: RELPAGE <= 12'd4095;
            12'd2484: RELPAGE <= 12'd4095;
            12'd2485: RELPAGE <= 12'd4095;
            12'd2486: RELPAGE <= 12'd4095;
            12'd2487: RELPAGE <= 12'd4095;
            12'd2488: RELPAGE <= 12'd4095;
            12'd2489: RELPAGE <= 12'd4095;
            12'd2490: RELPAGE <= 12'd4095;
            12'd2491: RELPAGE <= 12'd4095;
            12'd2492: RELPAGE <= 12'd4095;
            12'd2493: RELPAGE <= 12'd4095;
            12'd2494: RELPAGE <= 12'd4095;
            12'd2495: RELPAGE <= 12'd4095;
            12'd2496: RELPAGE <= 12'd4095;
            12'd2497: RELPAGE <= 12'd4095;
            12'd2498: RELPAGE <= 12'd4095;
            12'd2499: RELPAGE <= 12'd4095;
            12'd2500: RELPAGE <= 12'd4095;
            12'd2501: RELPAGE <= 12'd4095;
            12'd2502: RELPAGE <= 12'd4095;
            12'd2503: RELPAGE <= 12'd4095;
            12'd2504: RELPAGE <= 12'd4095;
            12'd2505: RELPAGE <= 12'd4095;
            12'd2506: RELPAGE <= 12'd4095;
            12'd2507: RELPAGE <= 12'd4095;
            12'd2508: RELPAGE <= 12'd4095;
            12'd2509: RELPAGE <= 12'd4095;
            12'd2510: RELPAGE <= 12'd4095;
            12'd2511: RELPAGE <= 12'd4095;
            12'd2512: RELPAGE <= 12'd4095;
            12'd2513: RELPAGE <= 12'd4095;
            12'd2514: RELPAGE <= 12'd4095;
            12'd2515: RELPAGE <= 12'd4095;
            12'd2516: RELPAGE <= 12'd4095;
            12'd2517: RELPAGE <= 12'd4095;
            12'd2518: RELPAGE <= 12'd4095;
            12'd2519: RELPAGE <= 12'd4095;
            12'd2520: RELPAGE <= 12'd4095;
            12'd2521: RELPAGE <= 12'd4095;
            12'd2522: RELPAGE <= 12'd4095;
            12'd2523: RELPAGE <= 12'd4095;
            12'd2524: RELPAGE <= 12'd4095;
            12'd2525: RELPAGE <= 12'd4095;
            12'd2526: RELPAGE <= 12'd4095;
            12'd2527: RELPAGE <= 12'd4095;
            12'd2528: RELPAGE <= 12'd4095;
            12'd2529: RELPAGE <= 12'd4095;
            12'd2530: RELPAGE <= 12'd4095;
            12'd2531: RELPAGE <= 12'd4095;
            12'd2532: RELPAGE <= 12'd4095;
            12'd2533: RELPAGE <= 12'd4095;
            12'd2534: RELPAGE <= 12'd4095;
            12'd2535: RELPAGE <= 12'd4095;
            12'd2536: RELPAGE <= 12'd4095;
            12'd2537: RELPAGE <= 12'd4095;
            12'd2538: RELPAGE <= 12'd4095;
            12'd2539: RELPAGE <= 12'd4095;
            12'd2540: RELPAGE <= 12'd4095;
            12'd2541: RELPAGE <= 12'd4095;
            12'd2542: RELPAGE <= 12'd4095;
            12'd2543: RELPAGE <= 12'd4095;
            12'd2544: RELPAGE <= 12'd4095;
            12'd2545: RELPAGE <= 12'd4095;
            12'd2546: RELPAGE <= 12'd4095;
            12'd2547: RELPAGE <= 12'd4095;
            12'd2548: RELPAGE <= 12'd4095;
            12'd2549: RELPAGE <= 12'd4095;
            12'd2550: RELPAGE <= 12'd4095;
            12'd2551: RELPAGE <= 12'd4095;
            12'd2552: RELPAGE <= 12'd4095;
            12'd2553: RELPAGE <= 12'd4095;
            12'd2554: RELPAGE <= 12'd4095;
            12'd2555: RELPAGE <= 12'd4095;
            12'd2556: RELPAGE <= 12'd4095;
            12'd2557: RELPAGE <= 12'd4095;
            12'd2558: RELPAGE <= 12'd4095;
            12'd2559: RELPAGE <= 12'd4095;
            12'd2560: RELPAGE <= 12'd4095;
            12'd2561: RELPAGE <= 12'd4095;
            12'd2562: RELPAGE <= 12'd4095;
            12'd2563: RELPAGE <= 12'd4095;
            12'd2564: RELPAGE <= 12'd4095;
            12'd2565: RELPAGE <= 12'd4095;
            12'd2566: RELPAGE <= 12'd4095;
            12'd2567: RELPAGE <= 12'd4095;
            12'd2568: RELPAGE <= 12'd4095;
            12'd2569: RELPAGE <= 12'd4095;
            12'd2570: RELPAGE <= 12'd4095;
            12'd2571: RELPAGE <= 12'd4095;
            12'd2572: RELPAGE <= 12'd4095;
            12'd2573: RELPAGE <= 12'd4095;
            12'd2574: RELPAGE <= 12'd4095;
            12'd2575: RELPAGE <= 12'd4095;
            12'd2576: RELPAGE <= 12'd4095;
            12'd2577: RELPAGE <= 12'd4095;
            12'd2578: RELPAGE <= 12'd4095;
            12'd2579: RELPAGE <= 12'd4095;
            12'd2580: RELPAGE <= 12'd4095;
            12'd2581: RELPAGE <= 12'd4095;
            12'd2582: RELPAGE <= 12'd4095;
            12'd2583: RELPAGE <= 12'd4095;
            12'd2584: RELPAGE <= 12'd4095;
            12'd2585: RELPAGE <= 12'd4095;
            12'd2586: RELPAGE <= 12'd4095;
            12'd2587: RELPAGE <= 12'd4095;
            12'd2588: RELPAGE <= 12'd4095;
            12'd2589: RELPAGE <= 12'd4095;
            12'd2590: RELPAGE <= 12'd4095;
            12'd2591: RELPAGE <= 12'd4095;
            12'd2592: RELPAGE <= 12'd4095;
            12'd2593: RELPAGE <= 12'd4095;
            12'd2594: RELPAGE <= 12'd4095;
            12'd2595: RELPAGE <= 12'd4095;
            12'd2596: RELPAGE <= 12'd4095;
            12'd2597: RELPAGE <= 12'd4095;
            12'd2598: RELPAGE <= 12'd4095;
            12'd2599: RELPAGE <= 12'd4095;
            12'd2600: RELPAGE <= 12'd4095;
            12'd2601: RELPAGE <= 12'd4095;
            12'd2602: RELPAGE <= 12'd4095;
            12'd2603: RELPAGE <= 12'd4095;
            12'd2604: RELPAGE <= 12'd4095;
            12'd2605: RELPAGE <= 12'd4095;
            12'd2606: RELPAGE <= 12'd4095;
            12'd2607: RELPAGE <= 12'd4095;
            12'd2608: RELPAGE <= 12'd4095;
            12'd2609: RELPAGE <= 12'd4095;
            12'd2610: RELPAGE <= 12'd4095;
            12'd2611: RELPAGE <= 12'd4095;
            12'd2612: RELPAGE <= 12'd4095;
            12'd2613: RELPAGE <= 12'd4095;
            12'd2614: RELPAGE <= 12'd4095;
            12'd2615: RELPAGE <= 12'd4095;
            12'd2616: RELPAGE <= 12'd4095;
            12'd2617: RELPAGE <= 12'd4095;
            12'd2618: RELPAGE <= 12'd4095;
            12'd2619: RELPAGE <= 12'd4095;
            12'd2620: RELPAGE <= 12'd4095;
            12'd2621: RELPAGE <= 12'd4095;
            12'd2622: RELPAGE <= 12'd4095;
            12'd2623: RELPAGE <= 12'd4095;
            12'd2624: RELPAGE <= 12'd4095;
            12'd2625: RELPAGE <= 12'd4095;
            12'd2626: RELPAGE <= 12'd4095;
            12'd2627: RELPAGE <= 12'd4095;
            12'd2628: RELPAGE <= 12'd4095;
            12'd2629: RELPAGE <= 12'd4095;
            12'd2630: RELPAGE <= 12'd4095;
            12'd2631: RELPAGE <= 12'd4095;
            12'd2632: RELPAGE <= 12'd4095;
            12'd2633: RELPAGE <= 12'd4095;
            12'd2634: RELPAGE <= 12'd4095;
            12'd2635: RELPAGE <= 12'd4095;
            12'd2636: RELPAGE <= 12'd4095;
            12'd2637: RELPAGE <= 12'd4095;
            12'd2638: RELPAGE <= 12'd4095;
            12'd2639: RELPAGE <= 12'd4095;
            12'd2640: RELPAGE <= 12'd4095;
            12'd2641: RELPAGE <= 12'd4095;
            12'd2642: RELPAGE <= 12'd4095;
            12'd2643: RELPAGE <= 12'd4095;
            12'd2644: RELPAGE <= 12'd4095;
            12'd2645: RELPAGE <= 12'd4095;
            12'd2646: RELPAGE <= 12'd4095;
            12'd2647: RELPAGE <= 12'd4095;
            12'd2648: RELPAGE <= 12'd4095;
            12'd2649: RELPAGE <= 12'd4095;
            12'd2650: RELPAGE <= 12'd4095;
            12'd2651: RELPAGE <= 12'd4095;
            12'd2652: RELPAGE <= 12'd4095;
            12'd2653: RELPAGE <= 12'd4095;
            12'd2654: RELPAGE <= 12'd4095;
            12'd2655: RELPAGE <= 12'd4095;
            12'd2656: RELPAGE <= 12'd4095;
            12'd2657: RELPAGE <= 12'd4095;
            12'd2658: RELPAGE <= 12'd4095;
            12'd2659: RELPAGE <= 12'd4095;
            12'd2660: RELPAGE <= 12'd4095;
            12'd2661: RELPAGE <= 12'd4095;
            12'd2662: RELPAGE <= 12'd4095;
            12'd2663: RELPAGE <= 12'd4095;
            12'd2664: RELPAGE <= 12'd4095;
            12'd2665: RELPAGE <= 12'd4095;
            12'd2666: RELPAGE <= 12'd4095;
            12'd2667: RELPAGE <= 12'd4095;
            12'd2668: RELPAGE <= 12'd4095;
            12'd2669: RELPAGE <= 12'd4095;
            12'd2670: RELPAGE <= 12'd4095;
            12'd2671: RELPAGE <= 12'd4095;
            12'd2672: RELPAGE <= 12'd4095;
            12'd2673: RELPAGE <= 12'd4095;
            12'd2674: RELPAGE <= 12'd4095;
            12'd2675: RELPAGE <= 12'd4095;
            12'd2676: RELPAGE <= 12'd4095;
            12'd2677: RELPAGE <= 12'd4095;
            12'd2678: RELPAGE <= 12'd4095;
            12'd2679: RELPAGE <= 12'd4095;
            12'd2680: RELPAGE <= 12'd4095;
            12'd2681: RELPAGE <= 12'd4095;
            12'd2682: RELPAGE <= 12'd4095;
            12'd2683: RELPAGE <= 12'd4095;
            12'd2684: RELPAGE <= 12'd4095;
            12'd2685: RELPAGE <= 12'd4095;
            12'd2686: RELPAGE <= 12'd4095;
            12'd2687: RELPAGE <= 12'd4095;
            12'd2688: RELPAGE <= 12'd4095;
            12'd2689: RELPAGE <= 12'd4095;
            12'd2690: RELPAGE <= 12'd4095;
            12'd2691: RELPAGE <= 12'd4095;
            12'd2692: RELPAGE <= 12'd4095;
            12'd2693: RELPAGE <= 12'd4095;
            12'd2694: RELPAGE <= 12'd4095;
            12'd2695: RELPAGE <= 12'd4095;
            12'd2696: RELPAGE <= 12'd4095;
            12'd2697: RELPAGE <= 12'd4095;
            12'd2698: RELPAGE <= 12'd4095;
            12'd2699: RELPAGE <= 12'd4095;
            12'd2700: RELPAGE <= 12'd4095;
            12'd2701: RELPAGE <= 12'd4095;
            12'd2702: RELPAGE <= 12'd4095;
            12'd2703: RELPAGE <= 12'd4095;
            12'd2704: RELPAGE <= 12'd4095;
            12'd2705: RELPAGE <= 12'd4095;
            12'd2706: RELPAGE <= 12'd4095;
            12'd2707: RELPAGE <= 12'd4095;
            12'd2708: RELPAGE <= 12'd4095;
            12'd2709: RELPAGE <= 12'd4095;
            12'd2710: RELPAGE <= 12'd4095;
            12'd2711: RELPAGE <= 12'd4095;
            12'd2712: RELPAGE <= 12'd4095;
            12'd2713: RELPAGE <= 12'd4095;
            12'd2714: RELPAGE <= 12'd4095;
            12'd2715: RELPAGE <= 12'd4095;
            12'd2716: RELPAGE <= 12'd4095;
            12'd2717: RELPAGE <= 12'd4095;
            12'd2718: RELPAGE <= 12'd4095;
            12'd2719: RELPAGE <= 12'd4095;
            12'd2720: RELPAGE <= 12'd4095;
            12'd2721: RELPAGE <= 12'd4095;
            12'd2722: RELPAGE <= 12'd4095;
            12'd2723: RELPAGE <= 12'd4095;
            12'd2724: RELPAGE <= 12'd4095;
            12'd2725: RELPAGE <= 12'd4095;
            12'd2726: RELPAGE <= 12'd4095;
            12'd2727: RELPAGE <= 12'd4095;
            12'd2728: RELPAGE <= 12'd4095;
            12'd2729: RELPAGE <= 12'd4095;
            12'd2730: RELPAGE <= 12'd4095;
            12'd2731: RELPAGE <= 12'd4095;
            12'd2732: RELPAGE <= 12'd4095;
            12'd2733: RELPAGE <= 12'd4095;
            12'd2734: RELPAGE <= 12'd4095;
            12'd2735: RELPAGE <= 12'd4095;
            12'd2736: RELPAGE <= 12'd4095;
            12'd2737: RELPAGE <= 12'd4095;
            12'd2738: RELPAGE <= 12'd4095;
            12'd2739: RELPAGE <= 12'd4095;
            12'd2740: RELPAGE <= 12'd4095;
            12'd2741: RELPAGE <= 12'd4095;
            12'd2742: RELPAGE <= 12'd4095;
            12'd2743: RELPAGE <= 12'd4095;
            12'd2744: RELPAGE <= 12'd4095;
            12'd2745: RELPAGE <= 12'd4095;
            12'd2746: RELPAGE <= 12'd4095;
            12'd2747: RELPAGE <= 12'd4095;
            12'd2748: RELPAGE <= 12'd4095;
            12'd2749: RELPAGE <= 12'd4095;
            12'd2750: RELPAGE <= 12'd4095;
            12'd2751: RELPAGE <= 12'd4095;
            12'd2752: RELPAGE <= 12'd4095;
            12'd2753: RELPAGE <= 12'd4095;
            12'd2754: RELPAGE <= 12'd4095;
            12'd2755: RELPAGE <= 12'd4095;
            12'd2756: RELPAGE <= 12'd4095;
            12'd2757: RELPAGE <= 12'd4095;
            12'd2758: RELPAGE <= 12'd4095;
            12'd2759: RELPAGE <= 12'd4095;
            12'd2760: RELPAGE <= 12'd4095;
            12'd2761: RELPAGE <= 12'd4095;
            12'd2762: RELPAGE <= 12'd4095;
            12'd2763: RELPAGE <= 12'd4095;
            12'd2764: RELPAGE <= 12'd4095;
            12'd2765: RELPAGE <= 12'd4095;
            12'd2766: RELPAGE <= 12'd4095;
            12'd2767: RELPAGE <= 12'd4095;
            12'd2768: RELPAGE <= 12'd4095;
            12'd2769: RELPAGE <= 12'd4095;
            12'd2770: RELPAGE <= 12'd4095;
            12'd2771: RELPAGE <= 12'd4095;
            12'd2772: RELPAGE <= 12'd4095;
            12'd2773: RELPAGE <= 12'd4095;
            12'd2774: RELPAGE <= 12'd4095;
            12'd2775: RELPAGE <= 12'd4095;
            12'd2776: RELPAGE <= 12'd4095;
            12'd2777: RELPAGE <= 12'd4095;
            12'd2778: RELPAGE <= 12'd4095;
            12'd2779: RELPAGE <= 12'd4095;
            12'd2780: RELPAGE <= 12'd4095;
            12'd2781: RELPAGE <= 12'd4095;
            12'd2782: RELPAGE <= 12'd4095;
            12'd2783: RELPAGE <= 12'd4095;
            12'd2784: RELPAGE <= 12'd4095;
            12'd2785: RELPAGE <= 12'd4095;
            12'd2786: RELPAGE <= 12'd4095;
            12'd2787: RELPAGE <= 12'd4095;
            12'd2788: RELPAGE <= 12'd4095;
            12'd2789: RELPAGE <= 12'd4095;
            12'd2790: RELPAGE <= 12'd4095;
            12'd2791: RELPAGE <= 12'd4095;
            12'd2792: RELPAGE <= 12'd4095;
            12'd2793: RELPAGE <= 12'd4095;
            12'd2794: RELPAGE <= 12'd4095;
            12'd2795: RELPAGE <= 12'd4095;
            12'd2796: RELPAGE <= 12'd4095;
            12'd2797: RELPAGE <= 12'd4095;
            12'd2798: RELPAGE <= 12'd4095;
            12'd2799: RELPAGE <= 12'd4095;
            12'd2800: RELPAGE <= 12'd4095;
            12'd2801: RELPAGE <= 12'd4095;
            12'd2802: RELPAGE <= 12'd4095;
            12'd2803: RELPAGE <= 12'd4095;
            12'd2804: RELPAGE <= 12'd4095;
            12'd2805: RELPAGE <= 12'd4095;
            12'd2806: RELPAGE <= 12'd4095;
            12'd2807: RELPAGE <= 12'd4095;
            12'd2808: RELPAGE <= 12'd4095;
            12'd2809: RELPAGE <= 12'd4095;
            12'd2810: RELPAGE <= 12'd4095;
            12'd2811: RELPAGE <= 12'd4095;
            12'd2812: RELPAGE <= 12'd4095;
            12'd2813: RELPAGE <= 12'd4095;
            12'd2814: RELPAGE <= 12'd4095;
            12'd2815: RELPAGE <= 12'd4095;
            12'd2816: RELPAGE <= 12'd4095;
            12'd2817: RELPAGE <= 12'd4095;
            12'd2818: RELPAGE <= 12'd4095;
            12'd2819: RELPAGE <= 12'd4095;
            12'd2820: RELPAGE <= 12'd4095;
            12'd2821: RELPAGE <= 12'd4095;
            12'd2822: RELPAGE <= 12'd4095;
            12'd2823: RELPAGE <= 12'd4095;
            12'd2824: RELPAGE <= 12'd4095;
            12'd2825: RELPAGE <= 12'd4095;
            12'd2826: RELPAGE <= 12'd4095;
            12'd2827: RELPAGE <= 12'd4095;
            12'd2828: RELPAGE <= 12'd4095;
            12'd2829: RELPAGE <= 12'd4095;
            12'd2830: RELPAGE <= 12'd4095;
            12'd2831: RELPAGE <= 12'd4095;
            12'd2832: RELPAGE <= 12'd4095;
            12'd2833: RELPAGE <= 12'd4095;
            12'd2834: RELPAGE <= 12'd4095;
            12'd2835: RELPAGE <= 12'd4095;
            12'd2836: RELPAGE <= 12'd4095;
            12'd2837: RELPAGE <= 12'd4095;
            12'd2838: RELPAGE <= 12'd4095;
            12'd2839: RELPAGE <= 12'd4095;
            12'd2840: RELPAGE <= 12'd4095;
            12'd2841: RELPAGE <= 12'd4095;
            12'd2842: RELPAGE <= 12'd4095;
            12'd2843: RELPAGE <= 12'd4095;
            12'd2844: RELPAGE <= 12'd4095;
            12'd2845: RELPAGE <= 12'd4095;
            12'd2846: RELPAGE <= 12'd4095;
            12'd2847: RELPAGE <= 12'd4095;
            12'd2848: RELPAGE <= 12'd4095;
            12'd2849: RELPAGE <= 12'd4095;
            12'd2850: RELPAGE <= 12'd4095;
            12'd2851: RELPAGE <= 12'd4095;
            12'd2852: RELPAGE <= 12'd4095;
            12'd2853: RELPAGE <= 12'd4095;
            12'd2854: RELPAGE <= 12'd4095;
            12'd2855: RELPAGE <= 12'd4095;
            12'd2856: RELPAGE <= 12'd4095;
            12'd2857: RELPAGE <= 12'd4095;
            12'd2858: RELPAGE <= 12'd4095;
            12'd2859: RELPAGE <= 12'd4095;
            12'd2860: RELPAGE <= 12'd4095;
            12'd2861: RELPAGE <= 12'd4095;
            12'd2862: RELPAGE <= 12'd4095;
            12'd2863: RELPAGE <= 12'd4095;
            12'd2864: RELPAGE <= 12'd4095;
            12'd2865: RELPAGE <= 12'd4095;
            12'd2866: RELPAGE <= 12'd4095;
            12'd2867: RELPAGE <= 12'd4095;
            12'd2868: RELPAGE <= 12'd4095;
            12'd2869: RELPAGE <= 12'd4095;
            12'd2870: RELPAGE <= 12'd4095;
            12'd2871: RELPAGE <= 12'd4095;
            12'd2872: RELPAGE <= 12'd4095;
            12'd2873: RELPAGE <= 12'd4095;
            12'd2874: RELPAGE <= 12'd4095;
            12'd2875: RELPAGE <= 12'd4095;
            12'd2876: RELPAGE <= 12'd4095;
            12'd2877: RELPAGE <= 12'd4095;
            12'd2878: RELPAGE <= 12'd4095;
            12'd2879: RELPAGE <= 12'd4095;
            12'd2880: RELPAGE <= 12'd4095;
            12'd2881: RELPAGE <= 12'd4095;
            12'd2882: RELPAGE <= 12'd4095;
            12'd2883: RELPAGE <= 12'd4095;
            12'd2884: RELPAGE <= 12'd4095;
            12'd2885: RELPAGE <= 12'd4095;
            12'd2886: RELPAGE <= 12'd4095;
            12'd2887: RELPAGE <= 12'd4095;
            12'd2888: RELPAGE <= 12'd4095;
            12'd2889: RELPAGE <= 12'd4095;
            12'd2890: RELPAGE <= 12'd4095;
            12'd2891: RELPAGE <= 12'd4095;
            12'd2892: RELPAGE <= 12'd4095;
            12'd2893: RELPAGE <= 12'd4095;
            12'd2894: RELPAGE <= 12'd4095;
            12'd2895: RELPAGE <= 12'd4095;
            12'd2896: RELPAGE <= 12'd4095;
            12'd2897: RELPAGE <= 12'd4095;
            12'd2898: RELPAGE <= 12'd4095;
            12'd2899: RELPAGE <= 12'd4095;
            12'd2900: RELPAGE <= 12'd4095;
            12'd2901: RELPAGE <= 12'd4095;
            12'd2902: RELPAGE <= 12'd4095;
            12'd2903: RELPAGE <= 12'd4095;
            12'd2904: RELPAGE <= 12'd4095;
            12'd2905: RELPAGE <= 12'd4095;
            12'd2906: RELPAGE <= 12'd4095;
            12'd2907: RELPAGE <= 12'd4095;
            12'd2908: RELPAGE <= 12'd4095;
            12'd2909: RELPAGE <= 12'd4095;
            12'd2910: RELPAGE <= 12'd4095;
            12'd2911: RELPAGE <= 12'd4095;
            12'd2912: RELPAGE <= 12'd4095;
            12'd2913: RELPAGE <= 12'd4095;
            12'd2914: RELPAGE <= 12'd4095;
            12'd2915: RELPAGE <= 12'd4095;
            12'd2916: RELPAGE <= 12'd4095;
            12'd2917: RELPAGE <= 12'd4095;
            12'd2918: RELPAGE <= 12'd4095;
            12'd2919: RELPAGE <= 12'd4095;
            12'd2920: RELPAGE <= 12'd4095;
            12'd2921: RELPAGE <= 12'd4095;
            12'd2922: RELPAGE <= 12'd4095;
            12'd2923: RELPAGE <= 12'd4095;
            12'd2924: RELPAGE <= 12'd4095;
            12'd2925: RELPAGE <= 12'd4095;
            12'd2926: RELPAGE <= 12'd4095;
            12'd2927: RELPAGE <= 12'd4095;
            12'd2928: RELPAGE <= 12'd4095;
            12'd2929: RELPAGE <= 12'd4095;
            12'd2930: RELPAGE <= 12'd4095;
            12'd2931: RELPAGE <= 12'd4095;
            12'd2932: RELPAGE <= 12'd4095;
            12'd2933: RELPAGE <= 12'd4095;
            12'd2934: RELPAGE <= 12'd4095;
            12'd2935: RELPAGE <= 12'd4095;
            12'd2936: RELPAGE <= 12'd4095;
            12'd2937: RELPAGE <= 12'd4095;
            12'd2938: RELPAGE <= 12'd4095;
            12'd2939: RELPAGE <= 12'd4095;
            12'd2940: RELPAGE <= 12'd4095;
            12'd2941: RELPAGE <= 12'd4095;
            12'd2942: RELPAGE <= 12'd4095;
            12'd2943: RELPAGE <= 12'd4095;
            12'd2944: RELPAGE <= 12'd4095;
            12'd2945: RELPAGE <= 12'd4095;
            12'd2946: RELPAGE <= 12'd4095;
            12'd2947: RELPAGE <= 12'd4095;
            12'd2948: RELPAGE <= 12'd4095;
            12'd2949: RELPAGE <= 12'd4095;
            12'd2950: RELPAGE <= 12'd4095;
            12'd2951: RELPAGE <= 12'd4095;
            12'd2952: RELPAGE <= 12'd4095;
            12'd2953: RELPAGE <= 12'd4095;
            12'd2954: RELPAGE <= 12'd4095;
            12'd2955: RELPAGE <= 12'd4095;
            12'd2956: RELPAGE <= 12'd4095;
            12'd2957: RELPAGE <= 12'd4095;
            12'd2958: RELPAGE <= 12'd4095;
            12'd2959: RELPAGE <= 12'd4095;
            12'd2960: RELPAGE <= 12'd4095;
            12'd2961: RELPAGE <= 12'd4095;
            12'd2962: RELPAGE <= 12'd4095;
            12'd2963: RELPAGE <= 12'd4095;
            12'd2964: RELPAGE <= 12'd4095;
            12'd2965: RELPAGE <= 12'd4095;
            12'd2966: RELPAGE <= 12'd4095;
            12'd2967: RELPAGE <= 12'd4095;
            12'd2968: RELPAGE <= 12'd4095;
            12'd2969: RELPAGE <= 12'd4095;
            12'd2970: RELPAGE <= 12'd4095;
            12'd2971: RELPAGE <= 12'd4095;
            12'd2972: RELPAGE <= 12'd4095;
            12'd2973: RELPAGE <= 12'd4095;
            12'd2974: RELPAGE <= 12'd4095;
            12'd2975: RELPAGE <= 12'd4095;
            12'd2976: RELPAGE <= 12'd4095;
            12'd2977: RELPAGE <= 12'd4095;
            12'd2978: RELPAGE <= 12'd4095;
            12'd2979: RELPAGE <= 12'd4095;
            12'd2980: RELPAGE <= 12'd4095;
            12'd2981: RELPAGE <= 12'd4095;
            12'd2982: RELPAGE <= 12'd4095;
            12'd2983: RELPAGE <= 12'd4095;
            12'd2984: RELPAGE <= 12'd4095;
            12'd2985: RELPAGE <= 12'd4095;
            12'd2986: RELPAGE <= 12'd4095;
            12'd2987: RELPAGE <= 12'd4095;
            12'd2988: RELPAGE <= 12'd4095;
            12'd2989: RELPAGE <= 12'd4095;
            12'd2990: RELPAGE <= 12'd4095;
            12'd2991: RELPAGE <= 12'd4095;
            12'd2992: RELPAGE <= 12'd4095;
            12'd2993: RELPAGE <= 12'd4095;
            12'd2994: RELPAGE <= 12'd4095;
            12'd2995: RELPAGE <= 12'd4095;
            12'd2996: RELPAGE <= 12'd4095;
            12'd2997: RELPAGE <= 12'd4095;
            12'd2998: RELPAGE <= 12'd4095;
            12'd2999: RELPAGE <= 12'd4095;
            12'd3000: RELPAGE <= 12'd4095;
            12'd3001: RELPAGE <= 12'd4095;
            12'd3002: RELPAGE <= 12'd4095;
            12'd3003: RELPAGE <= 12'd4095;
            12'd3004: RELPAGE <= 12'd4095;
            12'd3005: RELPAGE <= 12'd4095;
            12'd3006: RELPAGE <= 12'd4095;
            12'd3007: RELPAGE <= 12'd4095;
            12'd3008: RELPAGE <= 12'd4095;
            12'd3009: RELPAGE <= 12'd4095;
            12'd3010: RELPAGE <= 12'd4095;
            12'd3011: RELPAGE <= 12'd4095;
            12'd3012: RELPAGE <= 12'd4095;
            12'd3013: RELPAGE <= 12'd4095;
            12'd3014: RELPAGE <= 12'd4095;
            12'd3015: RELPAGE <= 12'd4095;
            12'd3016: RELPAGE <= 12'd4095;
            12'd3017: RELPAGE <= 12'd4095;
            12'd3018: RELPAGE <= 12'd4095;
            12'd3019: RELPAGE <= 12'd4095;
            12'd3020: RELPAGE <= 12'd4095;
            12'd3021: RELPAGE <= 12'd4095;
            12'd3022: RELPAGE <= 12'd4095;
            12'd3023: RELPAGE <= 12'd4095;
            12'd3024: RELPAGE <= 12'd4095;
            12'd3025: RELPAGE <= 12'd4095;
            12'd3026: RELPAGE <= 12'd4095;
            12'd3027: RELPAGE <= 12'd4095;
            12'd3028: RELPAGE <= 12'd4095;
            12'd3029: RELPAGE <= 12'd4095;
            12'd3030: RELPAGE <= 12'd4095;
            12'd3031: RELPAGE <= 12'd4095;
            12'd3032: RELPAGE <= 12'd4095;
            12'd3033: RELPAGE <= 12'd4095;
            12'd3034: RELPAGE <= 12'd4095;
            12'd3035: RELPAGE <= 12'd4095;
            12'd3036: RELPAGE <= 12'd4095;
            12'd3037: RELPAGE <= 12'd4095;
            12'd3038: RELPAGE <= 12'd4095;
            12'd3039: RELPAGE <= 12'd4095;
            12'd3040: RELPAGE <= 12'd4095;
            12'd3041: RELPAGE <= 12'd4095;
            12'd3042: RELPAGE <= 12'd4095;
            12'd3043: RELPAGE <= 12'd4095;
            12'd3044: RELPAGE <= 12'd4095;
            12'd3045: RELPAGE <= 12'd4095;
            12'd3046: RELPAGE <= 12'd4095;
            12'd3047: RELPAGE <= 12'd4095;
            12'd3048: RELPAGE <= 12'd4095;
            12'd3049: RELPAGE <= 12'd4095;
            12'd3050: RELPAGE <= 12'd4095;
            12'd3051: RELPAGE <= 12'd4095;
            12'd3052: RELPAGE <= 12'd4095;
            12'd3053: RELPAGE <= 12'd4095;
            12'd3054: RELPAGE <= 12'd4095;
            12'd3055: RELPAGE <= 12'd4095;
            12'd3056: RELPAGE <= 12'd4095;
            12'd3057: RELPAGE <= 12'd4095;
            12'd3058: RELPAGE <= 12'd4095;
            12'd3059: RELPAGE <= 12'd4095;
            12'd3060: RELPAGE <= 12'd4095;
            12'd3061: RELPAGE <= 12'd4095;
            12'd3062: RELPAGE <= 12'd4095;
            12'd3063: RELPAGE <= 12'd4095;
            12'd3064: RELPAGE <= 12'd4095;
            12'd3065: RELPAGE <= 12'd4095;
            12'd3066: RELPAGE <= 12'd4095;
            12'd3067: RELPAGE <= 12'd4095;
            12'd3068: RELPAGE <= 12'd4095;
            12'd3069: RELPAGE <= 12'd4095;
            12'd3070: RELPAGE <= 12'd4095;
            12'd3071: RELPAGE <= 12'd4095;
            12'd3072: RELPAGE <= 12'd4095;
            12'd3073: RELPAGE <= 12'd4095;
            12'd3074: RELPAGE <= 12'd4095;
            12'd3075: RELPAGE <= 12'd4095;
            12'd3076: RELPAGE <= 12'd4095;
            12'd3077: RELPAGE <= 12'd4095;
            12'd3078: RELPAGE <= 12'd4095;
            12'd3079: RELPAGE <= 12'd4095;
            12'd3080: RELPAGE <= 12'd4095;
            12'd3081: RELPAGE <= 12'd4095;
            12'd3082: RELPAGE <= 12'd4095;
            12'd3083: RELPAGE <= 12'd4095;
            12'd3084: RELPAGE <= 12'd4095;
            12'd3085: RELPAGE <= 12'd4095;
            12'd3086: RELPAGE <= 12'd4095;
            12'd3087: RELPAGE <= 12'd4095;
            12'd3088: RELPAGE <= 12'd4095;
            12'd3089: RELPAGE <= 12'd4095;
            12'd3090: RELPAGE <= 12'd4095;
            12'd3091: RELPAGE <= 12'd4095;
            12'd3092: RELPAGE <= 12'd4095;
            12'd3093: RELPAGE <= 12'd4095;
            12'd3094: RELPAGE <= 12'd4095;
            12'd3095: RELPAGE <= 12'd4095;
            12'd3096: RELPAGE <= 12'd4095;
            12'd3097: RELPAGE <= 12'd4095;
            12'd3098: RELPAGE <= 12'd4095;
            12'd3099: RELPAGE <= 12'd4095;
            12'd3100: RELPAGE <= 12'd4095;
            12'd3101: RELPAGE <= 12'd4095;
            12'd3102: RELPAGE <= 12'd4095;
            12'd3103: RELPAGE <= 12'd4095;
            12'd3104: RELPAGE <= 12'd4095;
            12'd3105: RELPAGE <= 12'd4095;
            12'd3106: RELPAGE <= 12'd4095;
            12'd3107: RELPAGE <= 12'd4095;
            12'd3108: RELPAGE <= 12'd4095;
            12'd3109: RELPAGE <= 12'd4095;
            12'd3110: RELPAGE <= 12'd4095;
            12'd3111: RELPAGE <= 12'd4095;
            12'd3112: RELPAGE <= 12'd4095;
            12'd3113: RELPAGE <= 12'd4095;
            12'd3114: RELPAGE <= 12'd4095;
            12'd3115: RELPAGE <= 12'd4095;
            12'd3116: RELPAGE <= 12'd4095;
            12'd3117: RELPAGE <= 12'd4095;
            12'd3118: RELPAGE <= 12'd4095;
            12'd3119: RELPAGE <= 12'd4095;
            12'd3120: RELPAGE <= 12'd4095;
            12'd3121: RELPAGE <= 12'd4095;
            12'd3122: RELPAGE <= 12'd4095;
            12'd3123: RELPAGE <= 12'd4095;
            12'd3124: RELPAGE <= 12'd4095;
            12'd3125: RELPAGE <= 12'd4095;
            12'd3126: RELPAGE <= 12'd4095;
            12'd3127: RELPAGE <= 12'd4095;
            12'd3128: RELPAGE <= 12'd4095;
            12'd3129: RELPAGE <= 12'd4095;
            12'd3130: RELPAGE <= 12'd4095;
            12'd3131: RELPAGE <= 12'd4095;
            12'd3132: RELPAGE <= 12'd4095;
            12'd3133: RELPAGE <= 12'd4095;
            12'd3134: RELPAGE <= 12'd4095;
            12'd3135: RELPAGE <= 12'd4095;
            12'd3136: RELPAGE <= 12'd4095;
            12'd3137: RELPAGE <= 12'd4095;
            12'd3138: RELPAGE <= 12'd4095;
            12'd3139: RELPAGE <= 12'd4095;
            12'd3140: RELPAGE <= 12'd4095;
            12'd3141: RELPAGE <= 12'd4095;
            12'd3142: RELPAGE <= 12'd4095;
            12'd3143: RELPAGE <= 12'd4095;
            12'd3144: RELPAGE <= 12'd4095;
            12'd3145: RELPAGE <= 12'd4095;
            12'd3146: RELPAGE <= 12'd4095;
            12'd3147: RELPAGE <= 12'd4095;
            12'd3148: RELPAGE <= 12'd4095;
            12'd3149: RELPAGE <= 12'd4095;
            12'd3150: RELPAGE <= 12'd4095;
            12'd3151: RELPAGE <= 12'd4095;
            12'd3152: RELPAGE <= 12'd4095;
            12'd3153: RELPAGE <= 12'd4095;
            12'd3154: RELPAGE <= 12'd4095;
            12'd3155: RELPAGE <= 12'd4095;
            12'd3156: RELPAGE <= 12'd4095;
            12'd3157: RELPAGE <= 12'd4095;
            12'd3158: RELPAGE <= 12'd4095;
            12'd3159: RELPAGE <= 12'd4095;
            12'd3160: RELPAGE <= 12'd4095;
            12'd3161: RELPAGE <= 12'd4095;
            12'd3162: RELPAGE <= 12'd4095;
            12'd3163: RELPAGE <= 12'd4095;
            12'd3164: RELPAGE <= 12'd4095;
            12'd3165: RELPAGE <= 12'd4095;
            12'd3166: RELPAGE <= 12'd4095;
            12'd3167: RELPAGE <= 12'd4095;
            12'd3168: RELPAGE <= 12'd4095;
            12'd3169: RELPAGE <= 12'd4095;
            12'd3170: RELPAGE <= 12'd4095;
            12'd3171: RELPAGE <= 12'd4095;
            12'd3172: RELPAGE <= 12'd4095;
            12'd3173: RELPAGE <= 12'd4095;
            12'd3174: RELPAGE <= 12'd4095;
            12'd3175: RELPAGE <= 12'd4095;
            12'd3176: RELPAGE <= 12'd4095;
            12'd3177: RELPAGE <= 12'd4095;
            12'd3178: RELPAGE <= 12'd4095;
            12'd3179: RELPAGE <= 12'd4095;
            12'd3180: RELPAGE <= 12'd4095;
            12'd3181: RELPAGE <= 12'd4095;
            12'd3182: RELPAGE <= 12'd4095;
            12'd3183: RELPAGE <= 12'd4095;
            12'd3184: RELPAGE <= 12'd4095;
            12'd3185: RELPAGE <= 12'd4095;
            12'd3186: RELPAGE <= 12'd4095;
            12'd3187: RELPAGE <= 12'd4095;
            12'd3188: RELPAGE <= 12'd4095;
            12'd3189: RELPAGE <= 12'd4095;
            12'd3190: RELPAGE <= 12'd4095;
            12'd3191: RELPAGE <= 12'd4095;
            12'd3192: RELPAGE <= 12'd4095;
            12'd3193: RELPAGE <= 12'd4095;
            12'd3194: RELPAGE <= 12'd4095;
            12'd3195: RELPAGE <= 12'd4095;
            12'd3196: RELPAGE <= 12'd4095;
            12'd3197: RELPAGE <= 12'd4095;
            12'd3198: RELPAGE <= 12'd4095;
            12'd3199: RELPAGE <= 12'd4095;
            12'd3200: RELPAGE <= 12'd4095;
            12'd3201: RELPAGE <= 12'd4095;
            12'd3202: RELPAGE <= 12'd4095;
            12'd3203: RELPAGE <= 12'd4095;
            12'd3204: RELPAGE <= 12'd4095;
            12'd3205: RELPAGE <= 12'd4095;
            12'd3206: RELPAGE <= 12'd4095;
            12'd3207: RELPAGE <= 12'd4095;
            12'd3208: RELPAGE <= 12'd4095;
            12'd3209: RELPAGE <= 12'd4095;
            12'd3210: RELPAGE <= 12'd4095;
            12'd3211: RELPAGE <= 12'd4095;
            12'd3212: RELPAGE <= 12'd4095;
            12'd3213: RELPAGE <= 12'd4095;
            12'd3214: RELPAGE <= 12'd4095;
            12'd3215: RELPAGE <= 12'd4095;
            12'd3216: RELPAGE <= 12'd4095;
            12'd3217: RELPAGE <= 12'd4095;
            12'd3218: RELPAGE <= 12'd4095;
            12'd3219: RELPAGE <= 12'd4095;
            12'd3220: RELPAGE <= 12'd4095;
            12'd3221: RELPAGE <= 12'd4095;
            12'd3222: RELPAGE <= 12'd4095;
            12'd3223: RELPAGE <= 12'd4095;
            12'd3224: RELPAGE <= 12'd4095;
            12'd3225: RELPAGE <= 12'd4095;
            12'd3226: RELPAGE <= 12'd4095;
            12'd3227: RELPAGE <= 12'd4095;
            12'd3228: RELPAGE <= 12'd4095;
            12'd3229: RELPAGE <= 12'd4095;
            12'd3230: RELPAGE <= 12'd4095;
            12'd3231: RELPAGE <= 12'd4095;
            12'd3232: RELPAGE <= 12'd4095;
            12'd3233: RELPAGE <= 12'd4095;
            12'd3234: RELPAGE <= 12'd4095;
            12'd3235: RELPAGE <= 12'd4095;
            12'd3236: RELPAGE <= 12'd4095;
            12'd3237: RELPAGE <= 12'd4095;
            12'd3238: RELPAGE <= 12'd4095;
            12'd3239: RELPAGE <= 12'd4095;
            12'd3240: RELPAGE <= 12'd4095;
            12'd3241: RELPAGE <= 12'd4095;
            12'd3242: RELPAGE <= 12'd4095;
            12'd3243: RELPAGE <= 12'd4095;
            12'd3244: RELPAGE <= 12'd4095;
            12'd3245: RELPAGE <= 12'd4095;
            12'd3246: RELPAGE <= 12'd4095;
            12'd3247: RELPAGE <= 12'd4095;
            12'd3248: RELPAGE <= 12'd4095;
            12'd3249: RELPAGE <= 12'd4095;
            12'd3250: RELPAGE <= 12'd4095;
            12'd3251: RELPAGE <= 12'd4095;
            12'd3252: RELPAGE <= 12'd4095;
            12'd3253: RELPAGE <= 12'd4095;
            12'd3254: RELPAGE <= 12'd4095;
            12'd3255: RELPAGE <= 12'd4095;
            12'd3256: RELPAGE <= 12'd4095;
            12'd3257: RELPAGE <= 12'd4095;
            12'd3258: RELPAGE <= 12'd4095;
            12'd3259: RELPAGE <= 12'd4095;
            12'd3260: RELPAGE <= 12'd4095;
            12'd3261: RELPAGE <= 12'd4095;
            12'd3262: RELPAGE <= 12'd4095;
            12'd3263: RELPAGE <= 12'd4095;
            12'd3264: RELPAGE <= 12'd4095;
            12'd3265: RELPAGE <= 12'd4095;
            12'd3266: RELPAGE <= 12'd4095;
            12'd3267: RELPAGE <= 12'd4095;
            12'd3268: RELPAGE <= 12'd4095;
            12'd3269: RELPAGE <= 12'd4095;
            12'd3270: RELPAGE <= 12'd4095;
            12'd3271: RELPAGE <= 12'd4095;
            12'd3272: RELPAGE <= 12'd4095;
            12'd3273: RELPAGE <= 12'd4095;
            12'd3274: RELPAGE <= 12'd4095;
            12'd3275: RELPAGE <= 12'd4095;
            12'd3276: RELPAGE <= 12'd4095;
            12'd3277: RELPAGE <= 12'd4095;
            12'd3278: RELPAGE <= 12'd4095;
            12'd3279: RELPAGE <= 12'd4095;
            12'd3280: RELPAGE <= 12'd4095;
            12'd3281: RELPAGE <= 12'd4095;
            12'd3282: RELPAGE <= 12'd4095;
            12'd3283: RELPAGE <= 12'd4095;
            12'd3284: RELPAGE <= 12'd4095;
            12'd3285: RELPAGE <= 12'd4095;
            12'd3286: RELPAGE <= 12'd4095;
            12'd3287: RELPAGE <= 12'd4095;
            12'd3288: RELPAGE <= 12'd4095;
            12'd3289: RELPAGE <= 12'd4095;
            12'd3290: RELPAGE <= 12'd4095;
            12'd3291: RELPAGE <= 12'd4095;
            12'd3292: RELPAGE <= 12'd4095;
            12'd3293: RELPAGE <= 12'd4095;
            12'd3294: RELPAGE <= 12'd4095;
            12'd3295: RELPAGE <= 12'd4095;
            12'd3296: RELPAGE <= 12'd4095;
            12'd3297: RELPAGE <= 12'd4095;
            12'd3298: RELPAGE <= 12'd4095;
            12'd3299: RELPAGE <= 12'd4095;
            12'd3300: RELPAGE <= 12'd4095;
            12'd3301: RELPAGE <= 12'd4095;
            12'd3302: RELPAGE <= 12'd4095;
            12'd3303: RELPAGE <= 12'd4095;
            12'd3304: RELPAGE <= 12'd4095;
            12'd3305: RELPAGE <= 12'd4095;
            12'd3306: RELPAGE <= 12'd4095;
            12'd3307: RELPAGE <= 12'd4095;
            12'd3308: RELPAGE <= 12'd4095;
            12'd3309: RELPAGE <= 12'd4095;
            12'd3310: RELPAGE <= 12'd4095;
            12'd3311: RELPAGE <= 12'd4095;
            12'd3312: RELPAGE <= 12'd4095;
            12'd3313: RELPAGE <= 12'd4095;
            12'd3314: RELPAGE <= 12'd4095;
            12'd3315: RELPAGE <= 12'd4095;
            12'd3316: RELPAGE <= 12'd4095;
            12'd3317: RELPAGE <= 12'd4095;
            12'd3318: RELPAGE <= 12'd4095;
            12'd3319: RELPAGE <= 12'd4095;
            12'd3320: RELPAGE <= 12'd4095;
            12'd3321: RELPAGE <= 12'd4095;
            12'd3322: RELPAGE <= 12'd4095;
            12'd3323: RELPAGE <= 12'd4095;
            12'd3324: RELPAGE <= 12'd4095;
            12'd3325: RELPAGE <= 12'd4095;
            12'd3326: RELPAGE <= 12'd4095;
            12'd3327: RELPAGE <= 12'd4095;
            12'd3328: RELPAGE <= 12'd4095;
            12'd3329: RELPAGE <= 12'd4095;
            12'd3330: RELPAGE <= 12'd4095;
            12'd3331: RELPAGE <= 12'd4095;
            12'd3332: RELPAGE <= 12'd4095;
            12'd3333: RELPAGE <= 12'd4095;
            12'd3334: RELPAGE <= 12'd4095;
            12'd3335: RELPAGE <= 12'd4095;
            12'd3336: RELPAGE <= 12'd4095;
            12'd3337: RELPAGE <= 12'd4095;
            12'd3338: RELPAGE <= 12'd4095;
            12'd3339: RELPAGE <= 12'd4095;
            12'd3340: RELPAGE <= 12'd4095;
            12'd3341: RELPAGE <= 12'd4095;
            12'd3342: RELPAGE <= 12'd4095;
            12'd3343: RELPAGE <= 12'd4095;
            12'd3344: RELPAGE <= 12'd4095;
            12'd3345: RELPAGE <= 12'd4095;
            12'd3346: RELPAGE <= 12'd4095;
            12'd3347: RELPAGE <= 12'd4095;
            12'd3348: RELPAGE <= 12'd4095;
            12'd3349: RELPAGE <= 12'd4095;
            12'd3350: RELPAGE <= 12'd4095;
            12'd3351: RELPAGE <= 12'd4095;
            12'd3352: RELPAGE <= 12'd4095;
            12'd3353: RELPAGE <= 12'd4095;
            12'd3354: RELPAGE <= 12'd4095;
            12'd3355: RELPAGE <= 12'd4095;
            12'd3356: RELPAGE <= 12'd4095;
            12'd3357: RELPAGE <= 12'd4095;
            12'd3358: RELPAGE <= 12'd4095;
            12'd3359: RELPAGE <= 12'd4095;
            12'd3360: RELPAGE <= 12'd4095;
            12'd3361: RELPAGE <= 12'd4095;
            12'd3362: RELPAGE <= 12'd4095;
            12'd3363: RELPAGE <= 12'd4095;
            12'd3364: RELPAGE <= 12'd4095;
            12'd3365: RELPAGE <= 12'd4095;
            12'd3366: RELPAGE <= 12'd4095;
            12'd3367: RELPAGE <= 12'd4095;
            12'd3368: RELPAGE <= 12'd4095;
            12'd3369: RELPAGE <= 12'd4095;
            12'd3370: RELPAGE <= 12'd4095;
            12'd3371: RELPAGE <= 12'd4095;
            12'd3372: RELPAGE <= 12'd4095;
            12'd3373: RELPAGE <= 12'd4095;
            12'd3374: RELPAGE <= 12'd4095;
            12'd3375: RELPAGE <= 12'd4095;
            12'd3376: RELPAGE <= 12'd4095;
            12'd3377: RELPAGE <= 12'd4095;
            12'd3378: RELPAGE <= 12'd4095;
            12'd3379: RELPAGE <= 12'd4095;
            12'd3380: RELPAGE <= 12'd4095;
            12'd3381: RELPAGE <= 12'd4095;
            12'd3382: RELPAGE <= 12'd4095;
            12'd3383: RELPAGE <= 12'd4095;
            12'd3384: RELPAGE <= 12'd4095;
            12'd3385: RELPAGE <= 12'd4095;
            12'd3386: RELPAGE <= 12'd4095;
            12'd3387: RELPAGE <= 12'd4095;
            12'd3388: RELPAGE <= 12'd4095;
            12'd3389: RELPAGE <= 12'd4095;
            12'd3390: RELPAGE <= 12'd4095;
            12'd3391: RELPAGE <= 12'd4095;
            12'd3392: RELPAGE <= 12'd4095;
            12'd3393: RELPAGE <= 12'd4095;
            12'd3394: RELPAGE <= 12'd4095;
            12'd3395: RELPAGE <= 12'd4095;
            12'd3396: RELPAGE <= 12'd4095;
            12'd3397: RELPAGE <= 12'd4095;
            12'd3398: RELPAGE <= 12'd4095;
            12'd3399: RELPAGE <= 12'd4095;
            12'd3400: RELPAGE <= 12'd4095;
            12'd3401: RELPAGE <= 12'd4095;
            12'd3402: RELPAGE <= 12'd4095;
            12'd3403: RELPAGE <= 12'd4095;
            12'd3404: RELPAGE <= 12'd4095;
            12'd3405: RELPAGE <= 12'd4095;
            12'd3406: RELPAGE <= 12'd4095;
            12'd3407: RELPAGE <= 12'd4095;
            12'd3408: RELPAGE <= 12'd4095;
            12'd3409: RELPAGE <= 12'd4095;
            12'd3410: RELPAGE <= 12'd4095;
            12'd3411: RELPAGE <= 12'd4095;
            12'd3412: RELPAGE <= 12'd4095;
            12'd3413: RELPAGE <= 12'd4095;
            12'd3414: RELPAGE <= 12'd4095;
            12'd3415: RELPAGE <= 12'd4095;
            12'd3416: RELPAGE <= 12'd4095;
            12'd3417: RELPAGE <= 12'd4095;
            12'd3418: RELPAGE <= 12'd4095;
            12'd3419: RELPAGE <= 12'd4095;
            12'd3420: RELPAGE <= 12'd4095;
            12'd3421: RELPAGE <= 12'd4095;
            12'd3422: RELPAGE <= 12'd4095;
            12'd3423: RELPAGE <= 12'd4095;
            12'd3424: RELPAGE <= 12'd4095;
            12'd3425: RELPAGE <= 12'd4095;
            12'd3426: RELPAGE <= 12'd4095;
            12'd3427: RELPAGE <= 12'd4095;
            12'd3428: RELPAGE <= 12'd4095;
            12'd3429: RELPAGE <= 12'd4095;
            12'd3430: RELPAGE <= 12'd4095;
            12'd3431: RELPAGE <= 12'd4095;
            12'd3432: RELPAGE <= 12'd4095;
            12'd3433: RELPAGE <= 12'd4095;
            12'd3434: RELPAGE <= 12'd4095;
            12'd3435: RELPAGE <= 12'd4095;
            12'd3436: RELPAGE <= 12'd4095;
            12'd3437: RELPAGE <= 12'd4095;
            12'd3438: RELPAGE <= 12'd4095;
            12'd3439: RELPAGE <= 12'd4095;
            12'd3440: RELPAGE <= 12'd4095;
            12'd3441: RELPAGE <= 12'd4095;
            12'd3442: RELPAGE <= 12'd4095;
            12'd3443: RELPAGE <= 12'd4095;
            12'd3444: RELPAGE <= 12'd4095;
            12'd3445: RELPAGE <= 12'd4095;
            12'd3446: RELPAGE <= 12'd4095;
            12'd3447: RELPAGE <= 12'd4095;
            12'd3448: RELPAGE <= 12'd4095;
            12'd3449: RELPAGE <= 12'd4095;
            12'd3450: RELPAGE <= 12'd4095;
            12'd3451: RELPAGE <= 12'd4095;
            12'd3452: RELPAGE <= 12'd4095;
            12'd3453: RELPAGE <= 12'd4095;
            12'd3454: RELPAGE <= 12'd4095;
            12'd3455: RELPAGE <= 12'd4095;
            12'd3456: RELPAGE <= 12'd4095;
            12'd3457: RELPAGE <= 12'd4095;
            12'd3458: RELPAGE <= 12'd4095;
            12'd3459: RELPAGE <= 12'd4095;
            12'd3460: RELPAGE <= 12'd4095;
            12'd3461: RELPAGE <= 12'd4095;
            12'd3462: RELPAGE <= 12'd4095;
            12'd3463: RELPAGE <= 12'd4095;
            12'd3464: RELPAGE <= 12'd4095;
            12'd3465: RELPAGE <= 12'd4095;
            12'd3466: RELPAGE <= 12'd4095;
            12'd3467: RELPAGE <= 12'd4095;
            12'd3468: RELPAGE <= 12'd4095;
            12'd3469: RELPAGE <= 12'd4095;
            12'd3470: RELPAGE <= 12'd4095;
            12'd3471: RELPAGE <= 12'd4095;
            12'd3472: RELPAGE <= 12'd4095;
            12'd3473: RELPAGE <= 12'd4095;
            12'd3474: RELPAGE <= 12'd4095;
            12'd3475: RELPAGE <= 12'd4095;
            12'd3476: RELPAGE <= 12'd4095;
            12'd3477: RELPAGE <= 12'd4095;
            12'd3478: RELPAGE <= 12'd4095;
            12'd3479: RELPAGE <= 12'd4095;
            12'd3480: RELPAGE <= 12'd4095;
            12'd3481: RELPAGE <= 12'd4095;
            12'd3482: RELPAGE <= 12'd4095;
            12'd3483: RELPAGE <= 12'd4095;
            12'd3484: RELPAGE <= 12'd4095;
            12'd3485: RELPAGE <= 12'd4095;
            12'd3486: RELPAGE <= 12'd4095;
            12'd3487: RELPAGE <= 12'd4095;
            12'd3488: RELPAGE <= 12'd4095;
            12'd3489: RELPAGE <= 12'd4095;
            12'd3490: RELPAGE <= 12'd4095;
            12'd3491: RELPAGE <= 12'd4095;
            12'd3492: RELPAGE <= 12'd4095;
            12'd3493: RELPAGE <= 12'd4095;
            12'd3494: RELPAGE <= 12'd4095;
            12'd3495: RELPAGE <= 12'd4095;
            12'd3496: RELPAGE <= 12'd4095;
            12'd3497: RELPAGE <= 12'd4095;
            12'd3498: RELPAGE <= 12'd4095;
            12'd3499: RELPAGE <= 12'd4095;
            12'd3500: RELPAGE <= 12'd4095;
            12'd3501: RELPAGE <= 12'd4095;
            12'd3502: RELPAGE <= 12'd4095;
            12'd3503: RELPAGE <= 12'd4095;
            12'd3504: RELPAGE <= 12'd4095;
            12'd3505: RELPAGE <= 12'd4095;
            12'd3506: RELPAGE <= 12'd4095;
            12'd3507: RELPAGE <= 12'd4095;
            12'd3508: RELPAGE <= 12'd4095;
            12'd3509: RELPAGE <= 12'd4095;
            12'd3510: RELPAGE <= 12'd4095;
            12'd3511: RELPAGE <= 12'd4095;
            12'd3512: RELPAGE <= 12'd4095;
            12'd3513: RELPAGE <= 12'd4095;
            12'd3514: RELPAGE <= 12'd4095;
            12'd3515: RELPAGE <= 12'd4095;
            12'd3516: RELPAGE <= 12'd4095;
            12'd3517: RELPAGE <= 12'd4095;
            12'd3518: RELPAGE <= 12'd4095;
            12'd3519: RELPAGE <= 12'd4095;
            12'd3520: RELPAGE <= 12'd4095;
            12'd3521: RELPAGE <= 12'd4095;
            12'd3522: RELPAGE <= 12'd4095;
            12'd3523: RELPAGE <= 12'd4095;
            12'd3524: RELPAGE <= 12'd4095;
            12'd3525: RELPAGE <= 12'd4095;
            12'd3526: RELPAGE <= 12'd4095;
            12'd3527: RELPAGE <= 12'd4095;
            12'd3528: RELPAGE <= 12'd4095;
            12'd3529: RELPAGE <= 12'd4095;
            12'd3530: RELPAGE <= 12'd4095;
            12'd3531: RELPAGE <= 12'd4095;
            12'd3532: RELPAGE <= 12'd4095;
            12'd3533: RELPAGE <= 12'd4095;
            12'd3534: RELPAGE <= 12'd4095;
            12'd3535: RELPAGE <= 12'd4095;
            12'd3536: RELPAGE <= 12'd4095;
            12'd3537: RELPAGE <= 12'd4095;
            12'd3538: RELPAGE <= 12'd4095;
            12'd3539: RELPAGE <= 12'd4095;
            12'd3540: RELPAGE <= 12'd4095;
            12'd3541: RELPAGE <= 12'd4095;
            12'd3542: RELPAGE <= 12'd4095;
            12'd3543: RELPAGE <= 12'd4095;
            12'd3544: RELPAGE <= 12'd4095;
            12'd3545: RELPAGE <= 12'd4095;
            12'd3546: RELPAGE <= 12'd4095;
            12'd3547: RELPAGE <= 12'd4095;
            12'd3548: RELPAGE <= 12'd4095;
            12'd3549: RELPAGE <= 12'd4095;
            12'd3550: RELPAGE <= 12'd4095;
            12'd3551: RELPAGE <= 12'd4095;
            12'd3552: RELPAGE <= 12'd4095;
            12'd3553: RELPAGE <= 12'd4095;
            12'd3554: RELPAGE <= 12'd4095;
            12'd3555: RELPAGE <= 12'd4095;
            12'd3556: RELPAGE <= 12'd4095;
            12'd3557: RELPAGE <= 12'd4095;
            12'd3558: RELPAGE <= 12'd4095;
            12'd3559: RELPAGE <= 12'd4095;
            12'd3560: RELPAGE <= 12'd4095;
            12'd3561: RELPAGE <= 12'd4095;
            12'd3562: RELPAGE <= 12'd4095;
            12'd3563: RELPAGE <= 12'd4095;
            12'd3564: RELPAGE <= 12'd4095;
            12'd3565: RELPAGE <= 12'd4095;
            12'd3566: RELPAGE <= 12'd4095;
            12'd3567: RELPAGE <= 12'd4095;
            12'd3568: RELPAGE <= 12'd4095;
            12'd3569: RELPAGE <= 12'd4095;
            12'd3570: RELPAGE <= 12'd4095;
            12'd3571: RELPAGE <= 12'd4095;
            12'd3572: RELPAGE <= 12'd4095;
            12'd3573: RELPAGE <= 12'd4095;
            12'd3574: RELPAGE <= 12'd4095;
            12'd3575: RELPAGE <= 12'd4095;
            12'd3576: RELPAGE <= 12'd4095;
            12'd3577: RELPAGE <= 12'd4095;
            12'd3578: RELPAGE <= 12'd4095;
            12'd3579: RELPAGE <= 12'd4095;
            12'd3580: RELPAGE <= 12'd4095;
            12'd3581: RELPAGE <= 12'd4095;
            12'd3582: RELPAGE <= 12'd4095;
            12'd3583: RELPAGE <= 12'd4095;
            12'd3584: RELPAGE <= 12'd4095;
            12'd3585: RELPAGE <= 12'd4095;
            12'd3586: RELPAGE <= 12'd4095;
            12'd3587: RELPAGE <= 12'd4095;
            12'd3588: RELPAGE <= 12'd4095;
            12'd3589: RELPAGE <= 12'd4095;
            12'd3590: RELPAGE <= 12'd4095;
            12'd3591: RELPAGE <= 12'd4095;
            12'd3592: RELPAGE <= 12'd4095;
            12'd3593: RELPAGE <= 12'd4095;
            12'd3594: RELPAGE <= 12'd4095;
            12'd3595: RELPAGE <= 12'd4095;
            12'd3596: RELPAGE <= 12'd4095;
            12'd3597: RELPAGE <= 12'd4095;
            12'd3598: RELPAGE <= 12'd4095;
            12'd3599: RELPAGE <= 12'd4095;
            12'd3600: RELPAGE <= 12'd4095;
            12'd3601: RELPAGE <= 12'd4095;
            12'd3602: RELPAGE <= 12'd4095;
            12'd3603: RELPAGE <= 12'd4095;
            12'd3604: RELPAGE <= 12'd4095;
            12'd3605: RELPAGE <= 12'd4095;
            12'd3606: RELPAGE <= 12'd4095;
            12'd3607: RELPAGE <= 12'd4095;
            12'd3608: RELPAGE <= 12'd4095;
            12'd3609: RELPAGE <= 12'd4095;
            12'd3610: RELPAGE <= 12'd4095;
            12'd3611: RELPAGE <= 12'd4095;
            12'd3612: RELPAGE <= 12'd4095;
            12'd3613: RELPAGE <= 12'd4095;
            12'd3614: RELPAGE <= 12'd4095;
            12'd3615: RELPAGE <= 12'd4095;
            12'd3616: RELPAGE <= 12'd4095;
            12'd3617: RELPAGE <= 12'd4095;
            12'd3618: RELPAGE <= 12'd4095;
            12'd3619: RELPAGE <= 12'd4095;
            12'd3620: RELPAGE <= 12'd4095;
            12'd3621: RELPAGE <= 12'd4095;
            12'd3622: RELPAGE <= 12'd4095;
            12'd3623: RELPAGE <= 12'd4095;
            12'd3624: RELPAGE <= 12'd4095;
            12'd3625: RELPAGE <= 12'd4095;
            12'd3626: RELPAGE <= 12'd4095;
            12'd3627: RELPAGE <= 12'd4095;
            12'd3628: RELPAGE <= 12'd4095;
            12'd3629: RELPAGE <= 12'd4095;
            12'd3630: RELPAGE <= 12'd4095;
            12'd3631: RELPAGE <= 12'd4095;
            12'd3632: RELPAGE <= 12'd4095;
            12'd3633: RELPAGE <= 12'd4095;
            12'd3634: RELPAGE <= 12'd4095;
            12'd3635: RELPAGE <= 12'd4095;
            12'd3636: RELPAGE <= 12'd4095;
            12'd3637: RELPAGE <= 12'd4095;
            12'd3638: RELPAGE <= 12'd4095;
            12'd3639: RELPAGE <= 12'd4095;
            12'd3640: RELPAGE <= 12'd4095;
            12'd3641: RELPAGE <= 12'd4095;
            12'd3642: RELPAGE <= 12'd4095;
            12'd3643: RELPAGE <= 12'd4095;
            12'd3644: RELPAGE <= 12'd4095;
            12'd3645: RELPAGE <= 12'd4095;
            12'd3646: RELPAGE <= 12'd4095;
            12'd3647: RELPAGE <= 12'd4095;
            12'd3648: RELPAGE <= 12'd4095;
            12'd3649: RELPAGE <= 12'd4095;
            12'd3650: RELPAGE <= 12'd4095;
            12'd3651: RELPAGE <= 12'd4095;
            12'd3652: RELPAGE <= 12'd4095;
            12'd3653: RELPAGE <= 12'd4095;
            12'd3654: RELPAGE <= 12'd4095;
            12'd3655: RELPAGE <= 12'd4095;
            12'd3656: RELPAGE <= 12'd4095;
            12'd3657: RELPAGE <= 12'd4095;
            12'd3658: RELPAGE <= 12'd4095;
            12'd3659: RELPAGE <= 12'd4095;
            12'd3660: RELPAGE <= 12'd4095;
            12'd3661: RELPAGE <= 12'd4095;
            12'd3662: RELPAGE <= 12'd4095;
            12'd3663: RELPAGE <= 12'd4095;
            12'd3664: RELPAGE <= 12'd4095;
            12'd3665: RELPAGE <= 12'd4095;
            12'd3666: RELPAGE <= 12'd4095;
            12'd3667: RELPAGE <= 12'd4095;
            12'd3668: RELPAGE <= 12'd4095;
            12'd3669: RELPAGE <= 12'd4095;
            12'd3670: RELPAGE <= 12'd4095;
            12'd3671: RELPAGE <= 12'd4095;
            12'd3672: RELPAGE <= 12'd4095;
            12'd3673: RELPAGE <= 12'd4095;
            12'd3674: RELPAGE <= 12'd4095;
            12'd3675: RELPAGE <= 12'd4095;
            12'd3676: RELPAGE <= 12'd4095;
            12'd3677: RELPAGE <= 12'd4095;
            12'd3678: RELPAGE <= 12'd4095;
            12'd3679: RELPAGE <= 12'd4095;
            12'd3680: RELPAGE <= 12'd4095;
            12'd3681: RELPAGE <= 12'd4095;
            12'd3682: RELPAGE <= 12'd4095;
            12'd3683: RELPAGE <= 12'd4095;
            12'd3684: RELPAGE <= 12'd4095;
            12'd3685: RELPAGE <= 12'd4095;
            12'd3686: RELPAGE <= 12'd4095;
            12'd3687: RELPAGE <= 12'd4095;
            12'd3688: RELPAGE <= 12'd4095;
            12'd3689: RELPAGE <= 12'd4095;
            12'd3690: RELPAGE <= 12'd4095;
            12'd3691: RELPAGE <= 12'd4095;
            12'd3692: RELPAGE <= 12'd4095;
            12'd3693: RELPAGE <= 12'd4095;
            12'd3694: RELPAGE <= 12'd4095;
            12'd3695: RELPAGE <= 12'd4095;
            12'd3696: RELPAGE <= 12'd4095;
            12'd3697: RELPAGE <= 12'd4095;
            12'd3698: RELPAGE <= 12'd4095;
            12'd3699: RELPAGE <= 12'd4095;
            12'd3700: RELPAGE <= 12'd4095;
            12'd3701: RELPAGE <= 12'd4095;
            12'd3702: RELPAGE <= 12'd4095;
            12'd3703: RELPAGE <= 12'd4095;
            12'd3704: RELPAGE <= 12'd4095;
            12'd3705: RELPAGE <= 12'd4095;
            12'd3706: RELPAGE <= 12'd4095;
            12'd3707: RELPAGE <= 12'd4095;
            12'd3708: RELPAGE <= 12'd4095;
            12'd3709: RELPAGE <= 12'd4095;
            12'd3710: RELPAGE <= 12'd4095;
            12'd3711: RELPAGE <= 12'd4095;
            12'd3712: RELPAGE <= 12'd4095;
            12'd3713: RELPAGE <= 12'd4095;
            12'd3714: RELPAGE <= 12'd4095;
            12'd3715: RELPAGE <= 12'd4095;
            12'd3716: RELPAGE <= 12'd4095;
            12'd3717: RELPAGE <= 12'd4095;
            12'd3718: RELPAGE <= 12'd4095;
            12'd3719: RELPAGE <= 12'd4095;
            12'd3720: RELPAGE <= 12'd4095;
            12'd3721: RELPAGE <= 12'd4095;
            12'd3722: RELPAGE <= 12'd4095;
            12'd3723: RELPAGE <= 12'd4095;
            12'd3724: RELPAGE <= 12'd4095;
            12'd3725: RELPAGE <= 12'd4095;
            12'd3726: RELPAGE <= 12'd4095;
            12'd3727: RELPAGE <= 12'd4095;
            12'd3728: RELPAGE <= 12'd4095;
            12'd3729: RELPAGE <= 12'd4095;
            12'd3730: RELPAGE <= 12'd4095;
            12'd3731: RELPAGE <= 12'd4095;
            12'd3732: RELPAGE <= 12'd4095;
            12'd3733: RELPAGE <= 12'd4095;
            12'd3734: RELPAGE <= 12'd4095;
            12'd3735: RELPAGE <= 12'd4095;
            12'd3736: RELPAGE <= 12'd4095;
            12'd3737: RELPAGE <= 12'd4095;
            12'd3738: RELPAGE <= 12'd4095;
            12'd3739: RELPAGE <= 12'd4095;
            12'd3740: RELPAGE <= 12'd4095;
            12'd3741: RELPAGE <= 12'd4095;
            12'd3742: RELPAGE <= 12'd4095;
            12'd3743: RELPAGE <= 12'd4095;
            12'd3744: RELPAGE <= 12'd4095;
            12'd3745: RELPAGE <= 12'd4095;
            12'd3746: RELPAGE <= 12'd4095;
            12'd3747: RELPAGE <= 12'd4095;
            12'd3748: RELPAGE <= 12'd4095;
            12'd3749: RELPAGE <= 12'd4095;
            12'd3750: RELPAGE <= 12'd4095;
            12'd3751: RELPAGE <= 12'd4095;
            12'd3752: RELPAGE <= 12'd4095;
            12'd3753: RELPAGE <= 12'd4095;
            12'd3754: RELPAGE <= 12'd4095;
            12'd3755: RELPAGE <= 12'd4095;
            12'd3756: RELPAGE <= 12'd4095;
            12'd3757: RELPAGE <= 12'd4095;
            12'd3758: RELPAGE <= 12'd4095;
            12'd3759: RELPAGE <= 12'd4095;
            12'd3760: RELPAGE <= 12'd4095;
            12'd3761: RELPAGE <= 12'd4095;
            12'd3762: RELPAGE <= 12'd4095;
            12'd3763: RELPAGE <= 12'd4095;
            12'd3764: RELPAGE <= 12'd4095;
            12'd3765: RELPAGE <= 12'd4095;
            12'd3766: RELPAGE <= 12'd4095;
            12'd3767: RELPAGE <= 12'd4095;
            12'd3768: RELPAGE <= 12'd4095;
            12'd3769: RELPAGE <= 12'd4095;
            12'd3770: RELPAGE <= 12'd4095;
            12'd3771: RELPAGE <= 12'd4095;
            12'd3772: RELPAGE <= 12'd4095;
            12'd3773: RELPAGE <= 12'd4095;
            12'd3774: RELPAGE <= 12'd4095;
            12'd3775: RELPAGE <= 12'd4095;
            12'd3776: RELPAGE <= 12'd4095;
            12'd3777: RELPAGE <= 12'd4095;
            12'd3778: RELPAGE <= 12'd4095;
            12'd3779: RELPAGE <= 12'd4095;
            12'd3780: RELPAGE <= 12'd4095;
            12'd3781: RELPAGE <= 12'd4095;
            12'd3782: RELPAGE <= 12'd4095;
            12'd3783: RELPAGE <= 12'd4095;
            12'd3784: RELPAGE <= 12'd4095;
            12'd3785: RELPAGE <= 12'd4095;
            12'd3786: RELPAGE <= 12'd4095;
            12'd3787: RELPAGE <= 12'd4095;
            12'd3788: RELPAGE <= 12'd4095;
            12'd3789: RELPAGE <= 12'd4095;
            12'd3790: RELPAGE <= 12'd4095;
            12'd3791: RELPAGE <= 12'd4095;
            12'd3792: RELPAGE <= 12'd4095;
            12'd3793: RELPAGE <= 12'd4095;
            12'd3794: RELPAGE <= 12'd4095;
            12'd3795: RELPAGE <= 12'd4095;
            12'd3796: RELPAGE <= 12'd4095;
            12'd3797: RELPAGE <= 12'd4095;
            12'd3798: RELPAGE <= 12'd4095;
            12'd3799: RELPAGE <= 12'd4095;
            12'd3800: RELPAGE <= 12'd4095;
            12'd3801: RELPAGE <= 12'd4095;
            12'd3802: RELPAGE <= 12'd4095;
            12'd3803: RELPAGE <= 12'd4095;
            12'd3804: RELPAGE <= 12'd4095;
            12'd3805: RELPAGE <= 12'd4095;
            12'd3806: RELPAGE <= 12'd4095;
            12'd3807: RELPAGE <= 12'd4095;
            12'd3808: RELPAGE <= 12'd4095;
            12'd3809: RELPAGE <= 12'd4095;
            12'd3810: RELPAGE <= 12'd4095;
            12'd3811: RELPAGE <= 12'd4095;
            12'd3812: RELPAGE <= 12'd4095;
            12'd3813: RELPAGE <= 12'd4095;
            12'd3814: RELPAGE <= 12'd4095;
            12'd3815: RELPAGE <= 12'd4095;
            12'd3816: RELPAGE <= 12'd4095;
            12'd3817: RELPAGE <= 12'd4095;
            12'd3818: RELPAGE <= 12'd4095;
            12'd3819: RELPAGE <= 12'd4095;
            12'd3820: RELPAGE <= 12'd4095;
            12'd3821: RELPAGE <= 12'd4095;
            12'd3822: RELPAGE <= 12'd4095;
            12'd3823: RELPAGE <= 12'd4095;
            12'd3824: RELPAGE <= 12'd4095;
            12'd3825: RELPAGE <= 12'd4095;
            12'd3826: RELPAGE <= 12'd4095;
            12'd3827: RELPAGE <= 12'd4095;
            12'd3828: RELPAGE <= 12'd4095;
            12'd3829: RELPAGE <= 12'd4095;
            12'd3830: RELPAGE <= 12'd4095;
            12'd3831: RELPAGE <= 12'd4095;
            12'd3832: RELPAGE <= 12'd4095;
            12'd3833: RELPAGE <= 12'd4095;
            12'd3834: RELPAGE <= 12'd4095;
            12'd3835: RELPAGE <= 12'd4095;
            12'd3836: RELPAGE <= 12'd4095;
            12'd3837: RELPAGE <= 12'd4095;
            12'd3838: RELPAGE <= 12'd4095;
            12'd3839: RELPAGE <= 12'd4095;
            12'd3840: RELPAGE <= 12'd4095;
            12'd3841: RELPAGE <= 12'd4095;
            12'd3842: RELPAGE <= 12'd4095;
            12'd3843: RELPAGE <= 12'd4095;
            12'd3844: RELPAGE <= 12'd4095;
            12'd3845: RELPAGE <= 12'd4095;
            12'd3846: RELPAGE <= 12'd4095;
            12'd3847: RELPAGE <= 12'd4095;
            12'd3848: RELPAGE <= 12'd4095;
            12'd3849: RELPAGE <= 12'd4095;
            12'd3850: RELPAGE <= 12'd4095;
            12'd3851: RELPAGE <= 12'd4095;
            12'd3852: RELPAGE <= 12'd4095;
            12'd3853: RELPAGE <= 12'd4095;
            12'd3854: RELPAGE <= 12'd4095;
            12'd3855: RELPAGE <= 12'd4095;
            12'd3856: RELPAGE <= 12'd4095;
            12'd3857: RELPAGE <= 12'd4095;
            12'd3858: RELPAGE <= 12'd4095;
            12'd3859: RELPAGE <= 12'd4095;
            12'd3860: RELPAGE <= 12'd4095;
            12'd3861: RELPAGE <= 12'd4095;
            12'd3862: RELPAGE <= 12'd4095;
            12'd3863: RELPAGE <= 12'd4095;
            12'd3864: RELPAGE <= 12'd4095;
            12'd3865: RELPAGE <= 12'd4095;
            12'd3866: RELPAGE <= 12'd4095;
            12'd3867: RELPAGE <= 12'd4095;
            12'd3868: RELPAGE <= 12'd4095;
            12'd3869: RELPAGE <= 12'd4095;
            12'd3870: RELPAGE <= 12'd4095;
            12'd3871: RELPAGE <= 12'd4095;
            12'd3872: RELPAGE <= 12'd4095;
            12'd3873: RELPAGE <= 12'd4095;
            12'd3874: RELPAGE <= 12'd4095;
            12'd3875: RELPAGE <= 12'd4095;
            12'd3876: RELPAGE <= 12'd4095;
            12'd3877: RELPAGE <= 12'd4095;
            12'd3878: RELPAGE <= 12'd4095;
            12'd3879: RELPAGE <= 12'd4095;
            12'd3880: RELPAGE <= 12'd4095;
            12'd3881: RELPAGE <= 12'd4095;
            12'd3882: RELPAGE <= 12'd4095;
            12'd3883: RELPAGE <= 12'd4095;
            12'd3884: RELPAGE <= 12'd4095;
            12'd3885: RELPAGE <= 12'd4095;
            12'd3886: RELPAGE <= 12'd4095;
            12'd3887: RELPAGE <= 12'd4095;
            12'd3888: RELPAGE <= 12'd4095;
            12'd3889: RELPAGE <= 12'd4095;
            12'd3890: RELPAGE <= 12'd4095;
            12'd3891: RELPAGE <= 12'd4095;
            12'd3892: RELPAGE <= 12'd4095;
            12'd3893: RELPAGE <= 12'd4095;
            12'd3894: RELPAGE <= 12'd4095;
            12'd3895: RELPAGE <= 12'd4095;
            12'd3896: RELPAGE <= 12'd4095;
            12'd3897: RELPAGE <= 12'd4095;
            12'd3898: RELPAGE <= 12'd4095;
            12'd3899: RELPAGE <= 12'd4095;
            12'd3900: RELPAGE <= 12'd4095;
            12'd3901: RELPAGE <= 12'd4095;
            12'd3902: RELPAGE <= 12'd4095;
            12'd3903: RELPAGE <= 12'd4095;
            12'd3904: RELPAGE <= 12'd4095;
            12'd3905: RELPAGE <= 12'd4095;
            12'd3906: RELPAGE <= 12'd4095;
            12'd3907: RELPAGE <= 12'd4095;
            12'd3908: RELPAGE <= 12'd4095;
            12'd3909: RELPAGE <= 12'd4095;
            12'd3910: RELPAGE <= 12'd4095;
            12'd3911: RELPAGE <= 12'd4095;
            12'd3912: RELPAGE <= 12'd4095;
            12'd3913: RELPAGE <= 12'd4095;
            12'd3914: RELPAGE <= 12'd4095;
            12'd3915: RELPAGE <= 12'd4095;
            12'd3916: RELPAGE <= 12'd4095;
            12'd3917: RELPAGE <= 12'd4095;
            12'd3918: RELPAGE <= 12'd4095;
            12'd3919: RELPAGE <= 12'd4095;
            12'd3920: RELPAGE <= 12'd4095;
            12'd3921: RELPAGE <= 12'd4095;
            12'd3922: RELPAGE <= 12'd4095;
            12'd3923: RELPAGE <= 12'd4095;
            12'd3924: RELPAGE <= 12'd4095;
            12'd3925: RELPAGE <= 12'd4095;
            12'd3926: RELPAGE <= 12'd4095;
            12'd3927: RELPAGE <= 12'd4095;
            12'd3928: RELPAGE <= 12'd4095;
            12'd3929: RELPAGE <= 12'd4095;
            12'd3930: RELPAGE <= 12'd4095;
            12'd3931: RELPAGE <= 12'd4095;
            12'd3932: RELPAGE <= 12'd4095;
            12'd3933: RELPAGE <= 12'd4095;
            12'd3934: RELPAGE <= 12'd4095;
            12'd3935: RELPAGE <= 12'd4095;
            12'd3936: RELPAGE <= 12'd4095;
            12'd3937: RELPAGE <= 12'd4095;
            12'd3938: RELPAGE <= 12'd4095;
            12'd3939: RELPAGE <= 12'd4095;
            12'd3940: RELPAGE <= 12'd4095;
            12'd3941: RELPAGE <= 12'd4095;
            12'd3942: RELPAGE <= 12'd4095;
            12'd3943: RELPAGE <= 12'd4095;
            12'd3944: RELPAGE <= 12'd4095;
            12'd3945: RELPAGE <= 12'd4095;
            12'd3946: RELPAGE <= 12'd4095;
            12'd3947: RELPAGE <= 12'd4095;
            12'd3948: RELPAGE <= 12'd4095;
            12'd3949: RELPAGE <= 12'd4095;
            12'd3950: RELPAGE <= 12'd4095;
            12'd3951: RELPAGE <= 12'd4095;
            12'd3952: RELPAGE <= 12'd4095;
            12'd3953: RELPAGE <= 12'd4095;
            12'd3954: RELPAGE <= 12'd4095;
            12'd3955: RELPAGE <= 12'd4095;
            12'd3956: RELPAGE <= 12'd4095;
            12'd3957: RELPAGE <= 12'd4095;
            12'd3958: RELPAGE <= 12'd4095;
            12'd3959: RELPAGE <= 12'd4095;
            12'd3960: RELPAGE <= 12'd4095;
            12'd3961: RELPAGE <= 12'd4095;
            12'd3962: RELPAGE <= 12'd4095;
            12'd3963: RELPAGE <= 12'd4095;
            12'd3964: RELPAGE <= 12'd4095;
            12'd3965: RELPAGE <= 12'd4095;
            12'd3966: RELPAGE <= 12'd4095;
            12'd3967: RELPAGE <= 12'd4095;
            12'd3968: RELPAGE <= 12'd4095;
            12'd3969: RELPAGE <= 12'd4095;
            12'd3970: RELPAGE <= 12'd4095;
            12'd3971: RELPAGE <= 12'd4095;
            12'd3972: RELPAGE <= 12'd4095;
            12'd3973: RELPAGE <= 12'd4095;
            12'd3974: RELPAGE <= 12'd4095;
            12'd3975: RELPAGE <= 12'd4095;
            12'd3976: RELPAGE <= 12'd4095;
            12'd3977: RELPAGE <= 12'd4095;
            12'd3978: RELPAGE <= 12'd4095;
            12'd3979: RELPAGE <= 12'd4095;
            12'd3980: RELPAGE <= 12'd4095;
            12'd3981: RELPAGE <= 12'd4095;
            12'd3982: RELPAGE <= 12'd4095;
            12'd3983: RELPAGE <= 12'd4095;
            12'd3984: RELPAGE <= 12'd4095;
            12'd3985: RELPAGE <= 12'd4095;
            12'd3986: RELPAGE <= 12'd4095;
            12'd3987: RELPAGE <= 12'd4095;
            12'd3988: RELPAGE <= 12'd4095;
            12'd3989: RELPAGE <= 12'd4095;
            12'd3990: RELPAGE <= 12'd4095;
            12'd3991: RELPAGE <= 12'd4095;
            12'd3992: RELPAGE <= 12'd4095;
            12'd3993: RELPAGE <= 12'd4095;
            12'd3994: RELPAGE <= 12'd4095;
            12'd3995: RELPAGE <= 12'd4095;
            12'd3996: RELPAGE <= 12'd4095;
            12'd3997: RELPAGE <= 12'd4095;
            12'd3998: RELPAGE <= 12'd4095;
            12'd3999: RELPAGE <= 12'd4095;
            12'd4000: RELPAGE <= 12'd4095;
            12'd4001: RELPAGE <= 12'd4095;
            12'd4002: RELPAGE <= 12'd4095;
            12'd4003: RELPAGE <= 12'd4095;
            12'd4004: RELPAGE <= 12'd4095;
            12'd4005: RELPAGE <= 12'd4095;
            12'd4006: RELPAGE <= 12'd4095;
            12'd4007: RELPAGE <= 12'd4095;
            12'd4008: RELPAGE <= 12'd4095;
            12'd4009: RELPAGE <= 12'd4095;
            12'd4010: RELPAGE <= 12'd4095;
            12'd4011: RELPAGE <= 12'd4095;
            12'd4012: RELPAGE <= 12'd4095;
            12'd4013: RELPAGE <= 12'd4095;
            12'd4014: RELPAGE <= 12'd4095;
            12'd4015: RELPAGE <= 12'd4095;
            12'd4016: RELPAGE <= 12'd4095;
            12'd4017: RELPAGE <= 12'd4095;
            12'd4018: RELPAGE <= 12'd4095;
            12'd4019: RELPAGE <= 12'd4095;
            12'd4020: RELPAGE <= 12'd4095;
            12'd4021: RELPAGE <= 12'd4095;
            12'd4022: RELPAGE <= 12'd4095;
            12'd4023: RELPAGE <= 12'd4095;
            12'd4024: RELPAGE <= 12'd4095;
            12'd4025: RELPAGE <= 12'd4095;
            12'd4026: RELPAGE <= 12'd4095;
            12'd4027: RELPAGE <= 12'd4095;
            12'd4028: RELPAGE <= 12'd4095;
            12'd4029: RELPAGE <= 12'd4095;
            12'd4030: RELPAGE <= 12'd4095;
            12'd4031: RELPAGE <= 12'd4095;
            12'd4032: RELPAGE <= 12'd4095;
            12'd4033: RELPAGE <= 12'd4095;
            12'd4034: RELPAGE <= 12'd4095;
            12'd4035: RELPAGE <= 12'd4095;
            12'd4036: RELPAGE <= 12'd4095;
            12'd4037: RELPAGE <= 12'd4095;
            12'd4038: RELPAGE <= 12'd4095;
            12'd4039: RELPAGE <= 12'd4095;
            12'd4040: RELPAGE <= 12'd4095;
            12'd4041: RELPAGE <= 12'd4095;
            12'd4042: RELPAGE <= 12'd4095;
            12'd4043: RELPAGE <= 12'd4095;
            12'd4044: RELPAGE <= 12'd4095;
            12'd4045: RELPAGE <= 12'd4095;
            12'd4046: RELPAGE <= 12'd4095;
            12'd4047: RELPAGE <= 12'd4095;
            12'd4048: RELPAGE <= 12'd4095;
            12'd4049: RELPAGE <= 12'd4095;
            12'd4050: RELPAGE <= 12'd4095;
            12'd4051: RELPAGE <= 12'd4095;
            12'd4052: RELPAGE <= 12'd4095;
            12'd4053: RELPAGE <= 12'd4095;
            12'd4054: RELPAGE <= 12'd4095;
            12'd4055: RELPAGE <= 12'd4095;
            12'd4056: RELPAGE <= 12'd4095;
            12'd4057: RELPAGE <= 12'd4095;
            12'd4058: RELPAGE <= 12'd4095;
            12'd4059: RELPAGE <= 12'd4095;
            12'd4060: RELPAGE <= 12'd4095;
            12'd4061: RELPAGE <= 12'd4095;
            12'd4062: RELPAGE <= 12'd4095;
            12'd4063: RELPAGE <= 12'd4095;
            12'd4064: RELPAGE <= 12'd4095;
            12'd4065: RELPAGE <= 12'd4095;
            12'd4066: RELPAGE <= 12'd4095;
            12'd4067: RELPAGE <= 12'd4095;
            12'd4068: RELPAGE <= 12'd4095;
            12'd4069: RELPAGE <= 12'd4095;
            12'd4070: RELPAGE <= 12'd4095;
            12'd4071: RELPAGE <= 12'd4095;
            12'd4072: RELPAGE <= 12'd4095;
            12'd4073: RELPAGE <= 12'd4095;
            12'd4074: RELPAGE <= 12'd4095;
            12'd4075: RELPAGE <= 12'd4095;
            12'd4076: RELPAGE <= 12'd4095;
            12'd4077: RELPAGE <= 12'd4095;
            12'd4078: RELPAGE <= 12'd4095;
            12'd4079: RELPAGE <= 12'd4095;
            12'd4080: RELPAGE <= 12'd4095;
            12'd4081: RELPAGE <= 12'd4095;
            12'd4082: RELPAGE <= 12'd4095;
            12'd4083: RELPAGE <= 12'd4095;
            12'd4084: RELPAGE <= 12'd4095;
            12'd4085: RELPAGE <= 12'd4095;
            12'd4086: RELPAGE <= 12'd4095;
            12'd4087: RELPAGE <= 12'd4095;
            12'd4088: RELPAGE <= 12'd4095;
            12'd4089: RELPAGE <= 12'd4095;
            12'd4090: RELPAGE <= 12'd4095;
            12'd4091: RELPAGE <= 12'd4095;
            12'd4092: RELPAGE <= 12'd4095;
            12'd4093: RELPAGE <= 12'd4095;
            12'd4094: RELPAGE <= 12'd4095;
            12'd4095: RELPAGE <= 12'd4095;
        endcase
    end
end

endmodule