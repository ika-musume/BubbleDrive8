module PositionPageConverter 
(
    input   wire            position_convert,
    input   wire    [11:0]  current_position,
    output  reg     [11:0]  current_page = 12'd4095
);

    always @ (posedge position_convert)
    begin
        case (current_position)
            12'd0: current_page <= 12'd1862;
            12'd1: current_page <= 12'd331;
            12'd2: current_page <= 12'd853;
            12'd3: current_page <= 12'd1375;
            12'd4: current_page <= 12'd1897;
            12'd5: current_page <= 12'd366;
            12'd6: current_page <= 12'd888;
            12'd7: current_page <= 12'd1410;
            12'd8: current_page <= 12'd1932;
            12'd9: current_page <= 12'd401;
            12'd10: current_page <= 12'd923;
            12'd11: current_page <= 12'd1445;
            12'd12: current_page <= 12'd1967;
            12'd13: current_page <= 12'd436;
            12'd14: current_page <= 12'd958;
            12'd15: current_page <= 12'd1480;
            12'd16: current_page <= 12'd2002;
            12'd17: current_page <= 12'd471;
            12'd18: current_page <= 12'd993;
            12'd19: current_page <= 12'd1515;
            12'd20: current_page <= 12'd2037;
            12'd21: current_page <= 12'd506;
            12'd22: current_page <= 12'd1028;
            12'd23: current_page <= 12'd1550;
            12'd24: current_page <= 12'd19;
            12'd25: current_page <= 12'd541;
            12'd26: current_page <= 12'd1063;
            12'd27: current_page <= 12'd1585;
            12'd28: current_page <= 12'd54;
            12'd29: current_page <= 12'd576;
            12'd30: current_page <= 12'd1098;
            12'd31: current_page <= 12'd1620;
            12'd32: current_page <= 12'd89;
            12'd33: current_page <= 12'd611;
            12'd34: current_page <= 12'd1133;
            12'd35: current_page <= 12'd1655;
            12'd36: current_page <= 12'd124;
            12'd37: current_page <= 12'd646;
            12'd38: current_page <= 12'd1168;
            12'd39: current_page <= 12'd1690;
            12'd40: current_page <= 12'd159;
            12'd41: current_page <= 12'd681;
            12'd42: current_page <= 12'd1203;
            12'd43: current_page <= 12'd1725;
            12'd44: current_page <= 12'd194;
            12'd45: current_page <= 12'd716;
            12'd46: current_page <= 12'd1238;
            12'd47: current_page <= 12'd1760;
            12'd48: current_page <= 12'd229;
            12'd49: current_page <= 12'd751;
            12'd50: current_page <= 12'd1273;
            12'd51: current_page <= 12'd1795;
            12'd52: current_page <= 12'd264;
            12'd53: current_page <= 12'd786;
            12'd54: current_page <= 12'd1308;
            12'd55: current_page <= 12'd1830;
            12'd56: current_page <= 12'd299;
            12'd57: current_page <= 12'd821;
            12'd58: current_page <= 12'd1343;
            12'd59: current_page <= 12'd1865;
            12'd60: current_page <= 12'd334;
            12'd61: current_page <= 12'd856;
            12'd62: current_page <= 12'd1378;
            12'd63: current_page <= 12'd1900;
            12'd64: current_page <= 12'd369;
            12'd65: current_page <= 12'd891;
            12'd66: current_page <= 12'd1413;
            12'd67: current_page <= 12'd1935;
            12'd68: current_page <= 12'd404;
            12'd69: current_page <= 12'd926;
            12'd70: current_page <= 12'd1448;
            12'd71: current_page <= 12'd1970;
            12'd72: current_page <= 12'd439;
            12'd73: current_page <= 12'd961;
            12'd74: current_page <= 12'd1483;
            12'd75: current_page <= 12'd2005;
            12'd76: current_page <= 12'd474;
            12'd77: current_page <= 12'd996;
            12'd78: current_page <= 12'd1518;
            12'd79: current_page <= 12'd2040;
            12'd80: current_page <= 12'd509;
            12'd81: current_page <= 12'd1031;
            12'd82: current_page <= 12'd1553;
            12'd83: current_page <= 12'd22;
            12'd84: current_page <= 12'd544;
            12'd85: current_page <= 12'd1066;
            12'd86: current_page <= 12'd1588;
            12'd87: current_page <= 12'd57;
            12'd88: current_page <= 12'd579;
            12'd89: current_page <= 12'd1101;
            12'd90: current_page <= 12'd1623;
            12'd91: current_page <= 12'd92;
            12'd92: current_page <= 12'd614;
            12'd93: current_page <= 12'd1136;
            12'd94: current_page <= 12'd1658;
            12'd95: current_page <= 12'd127;
            12'd96: current_page <= 12'd649;
            12'd97: current_page <= 12'd1171;
            12'd98: current_page <= 12'd1693;
            12'd99: current_page <= 12'd162;
            12'd100: current_page <= 12'd684;
            12'd101: current_page <= 12'd1206;
            12'd102: current_page <= 12'd1728;
            12'd103: current_page <= 12'd197;
            12'd104: current_page <= 12'd719;
            12'd105: current_page <= 12'd1241;
            12'd106: current_page <= 12'd1763;
            12'd107: current_page <= 12'd232;
            12'd108: current_page <= 12'd754;
            12'd109: current_page <= 12'd1276;
            12'd110: current_page <= 12'd1798;
            12'd111: current_page <= 12'd267;
            12'd112: current_page <= 12'd789;
            12'd113: current_page <= 12'd1311;
            12'd114: current_page <= 12'd1833;
            12'd115: current_page <= 12'd302;
            12'd116: current_page <= 12'd824;
            12'd117: current_page <= 12'd1346;
            12'd118: current_page <= 12'd1868;
            12'd119: current_page <= 12'd337;
            12'd120: current_page <= 12'd859;
            12'd121: current_page <= 12'd1381;
            12'd122: current_page <= 12'd1903;
            12'd123: current_page <= 12'd372;
            12'd124: current_page <= 12'd894;
            12'd125: current_page <= 12'd1416;
            12'd126: current_page <= 12'd1938;
            12'd127: current_page <= 12'd407;
            12'd128: current_page <= 12'd929;
            12'd129: current_page <= 12'd1451;
            12'd130: current_page <= 12'd1973;
            12'd131: current_page <= 12'd442;
            12'd132: current_page <= 12'd964;
            12'd133: current_page <= 12'd1486;
            12'd134: current_page <= 12'd2008;
            12'd135: current_page <= 12'd477;
            12'd136: current_page <= 12'd999;
            12'd137: current_page <= 12'd1521;
            12'd138: current_page <= 12'd2043;
            12'd139: current_page <= 12'd512;
            12'd140: current_page <= 12'd1034;
            12'd141: current_page <= 12'd1556;
            12'd142: current_page <= 12'd25;
            12'd143: current_page <= 12'd547;
            12'd144: current_page <= 12'd1069;
            12'd145: current_page <= 12'd1591;
            12'd146: current_page <= 12'd60;
            12'd147: current_page <= 12'd582;
            12'd148: current_page <= 12'd1104;
            12'd149: current_page <= 12'd1626;
            12'd150: current_page <= 12'd95;
            12'd151: current_page <= 12'd617;
            12'd152: current_page <= 12'd1139;
            12'd153: current_page <= 12'd1661;
            12'd154: current_page <= 12'd130;
            12'd155: current_page <= 12'd652;
            12'd156: current_page <= 12'd1174;
            12'd157: current_page <= 12'd1696;
            12'd158: current_page <= 12'd165;
            12'd159: current_page <= 12'd687;
            12'd160: current_page <= 12'd1209;
            12'd161: current_page <= 12'd1731;
            12'd162: current_page <= 12'd200;
            12'd163: current_page <= 12'd722;
            12'd164: current_page <= 12'd1244;
            12'd165: current_page <= 12'd1766;
            12'd166: current_page <= 12'd235;
            12'd167: current_page <= 12'd757;
            12'd168: current_page <= 12'd1279;
            12'd169: current_page <= 12'd1801;
            12'd170: current_page <= 12'd270;
            12'd171: current_page <= 12'd792;
            12'd172: current_page <= 12'd1314;
            12'd173: current_page <= 12'd1836;
            12'd174: current_page <= 12'd305;
            12'd175: current_page <= 12'd827;
            12'd176: current_page <= 12'd1349;
            12'd177: current_page <= 12'd1871;
            12'd178: current_page <= 12'd340;
            12'd179: current_page <= 12'd862;
            12'd180: current_page <= 12'd1384;
            12'd181: current_page <= 12'd1906;
            12'd182: current_page <= 12'd375;
            12'd183: current_page <= 12'd897;
            12'd184: current_page <= 12'd1419;
            12'd185: current_page <= 12'd1941;
            12'd186: current_page <= 12'd410;
            12'd187: current_page <= 12'd932;
            12'd188: current_page <= 12'd1454;
            12'd189: current_page <= 12'd1976;
            12'd190: current_page <= 12'd445;
            12'd191: current_page <= 12'd967;
            12'd192: current_page <= 12'd1489;
            12'd193: current_page <= 12'd2011;
            12'd194: current_page <= 12'd480;
            12'd195: current_page <= 12'd1002;
            12'd196: current_page <= 12'd1524;
            12'd197: current_page <= 12'd2046;
            12'd198: current_page <= 12'd515;
            12'd199: current_page <= 12'd1037;
            12'd200: current_page <= 12'd1559;
            12'd201: current_page <= 12'd28;
            12'd202: current_page <= 12'd550;
            12'd203: current_page <= 12'd1072;
            12'd204: current_page <= 12'd1594;
            12'd205: current_page <= 12'd63;
            12'd206: current_page <= 12'd585;
            12'd207: current_page <= 12'd1107;
            12'd208: current_page <= 12'd1629;
            12'd209: current_page <= 12'd98;
            12'd210: current_page <= 12'd620;
            12'd211: current_page <= 12'd1142;
            12'd212: current_page <= 12'd1664;
            12'd213: current_page <= 12'd133;
            12'd214: current_page <= 12'd655;
            12'd215: current_page <= 12'd1177;
            12'd216: current_page <= 12'd1699;
            12'd217: current_page <= 12'd168;
            12'd218: current_page <= 12'd690;
            12'd219: current_page <= 12'd1212;
            12'd220: current_page <= 12'd1734;
            12'd221: current_page <= 12'd203;
            12'd222: current_page <= 12'd725;
            12'd223: current_page <= 12'd1247;
            12'd224: current_page <= 12'd1769;
            12'd225: current_page <= 12'd238;
            12'd226: current_page <= 12'd760;
            12'd227: current_page <= 12'd1282;
            12'd228: current_page <= 12'd1804;
            12'd229: current_page <= 12'd273;
            12'd230: current_page <= 12'd795;
            12'd231: current_page <= 12'd1317;
            12'd232: current_page <= 12'd1839;
            12'd233: current_page <= 12'd308;
            12'd234: current_page <= 12'd830;
            12'd235: current_page <= 12'd1352;
            12'd236: current_page <= 12'd1874;
            12'd237: current_page <= 12'd343;
            12'd238: current_page <= 12'd865;
            12'd239: current_page <= 12'd1387;
            12'd240: current_page <= 12'd1909;
            12'd241: current_page <= 12'd378;
            12'd242: current_page <= 12'd900;
            12'd243: current_page <= 12'd1422;
            12'd244: current_page <= 12'd1944;
            12'd245: current_page <= 12'd413;
            12'd246: current_page <= 12'd935;
            12'd247: current_page <= 12'd1457;
            12'd248: current_page <= 12'd1979;
            12'd249: current_page <= 12'd448;
            12'd250: current_page <= 12'd970;
            12'd251: current_page <= 12'd1492;
            12'd252: current_page <= 12'd2014;
            12'd253: current_page <= 12'd483;
            12'd254: current_page <= 12'd1005;
            12'd255: current_page <= 12'd1527;
            12'd256: current_page <= 12'd2049;
            12'd257: current_page <= 12'd518;
            12'd258: current_page <= 12'd1040;
            12'd259: current_page <= 12'd1562;
            12'd260: current_page <= 12'd31;
            12'd261: current_page <= 12'd553;
            12'd262: current_page <= 12'd1075;
            12'd263: current_page <= 12'd1597;
            12'd264: current_page <= 12'd66;
            12'd265: current_page <= 12'd588;
            12'd266: current_page <= 12'd1110;
            12'd267: current_page <= 12'd1632;
            12'd268: current_page <= 12'd101;
            12'd269: current_page <= 12'd623;
            12'd270: current_page <= 12'd1145;
            12'd271: current_page <= 12'd1667;
            12'd272: current_page <= 12'd136;
            12'd273: current_page <= 12'd658;
            12'd274: current_page <= 12'd1180;
            12'd275: current_page <= 12'd1702;
            12'd276: current_page <= 12'd171;
            12'd277: current_page <= 12'd693;
            12'd278: current_page <= 12'd1215;
            12'd279: current_page <= 12'd1737;
            12'd280: current_page <= 12'd206;
            12'd281: current_page <= 12'd728;
            12'd282: current_page <= 12'd1250;
            12'd283: current_page <= 12'd1772;
            12'd284: current_page <= 12'd241;
            12'd285: current_page <= 12'd763;
            12'd286: current_page <= 12'd1285;
            12'd287: current_page <= 12'd1807;
            12'd288: current_page <= 12'd276;
            12'd289: current_page <= 12'd798;
            12'd290: current_page <= 12'd1320;
            12'd291: current_page <= 12'd1842;
            12'd292: current_page <= 12'd311;
            12'd293: current_page <= 12'd833;
            12'd294: current_page <= 12'd1355;
            12'd295: current_page <= 12'd1877;
            12'd296: current_page <= 12'd346;
            12'd297: current_page <= 12'd868;
            12'd298: current_page <= 12'd1390;
            12'd299: current_page <= 12'd1912;
            12'd300: current_page <= 12'd381;
            12'd301: current_page <= 12'd903;
            12'd302: current_page <= 12'd1425;
            12'd303: current_page <= 12'd1947;
            12'd304: current_page <= 12'd416;
            12'd305: current_page <= 12'd938;
            12'd306: current_page <= 12'd1460;
            12'd307: current_page <= 12'd1982;
            12'd308: current_page <= 12'd451;
            12'd309: current_page <= 12'd973;
            12'd310: current_page <= 12'd1495;
            12'd311: current_page <= 12'd2017;
            12'd312: current_page <= 12'd486;
            12'd313: current_page <= 12'd1008;
            12'd314: current_page <= 12'd1530;
            12'd315: current_page <= 12'd2052;
            12'd316: current_page <= 12'd521;
            12'd317: current_page <= 12'd1043;
            12'd318: current_page <= 12'd1565;
            12'd319: current_page <= 12'd34;
            12'd320: current_page <= 12'd556;
            12'd321: current_page <= 12'd1078;
            12'd322: current_page <= 12'd1600;
            12'd323: current_page <= 12'd69;
            12'd324: current_page <= 12'd591;
            12'd325: current_page <= 12'd1113;
            12'd326: current_page <= 12'd1635;
            12'd327: current_page <= 12'd104;
            12'd328: current_page <= 12'd626;
            12'd329: current_page <= 12'd1148;
            12'd330: current_page <= 12'd1670;
            12'd331: current_page <= 12'd139;
            12'd332: current_page <= 12'd661;
            12'd333: current_page <= 12'd1183;
            12'd334: current_page <= 12'd1705;
            12'd335: current_page <= 12'd174;
            12'd336: current_page <= 12'd696;
            12'd337: current_page <= 12'd1218;
            12'd338: current_page <= 12'd1740;
            12'd339: current_page <= 12'd209;
            12'd340: current_page <= 12'd731;
            12'd341: current_page <= 12'd1253;
            12'd342: current_page <= 12'd1775;
            12'd343: current_page <= 12'd244;
            12'd344: current_page <= 12'd766;
            12'd345: current_page <= 12'd1288;
            12'd346: current_page <= 12'd1810;
            12'd347: current_page <= 12'd279;
            12'd348: current_page <= 12'd801;
            12'd349: current_page <= 12'd1323;
            12'd350: current_page <= 12'd1845;
            12'd351: current_page <= 12'd314;
            12'd352: current_page <= 12'd836;
            12'd353: current_page <= 12'd1358;
            12'd354: current_page <= 12'd1880;
            12'd355: current_page <= 12'd349;
            12'd356: current_page <= 12'd871;
            12'd357: current_page <= 12'd1393;
            12'd358: current_page <= 12'd1915;
            12'd359: current_page <= 12'd384;
            12'd360: current_page <= 12'd906;
            12'd361: current_page <= 12'd1428;
            12'd362: current_page <= 12'd1950;
            12'd363: current_page <= 12'd419;
            12'd364: current_page <= 12'd941;
            12'd365: current_page <= 12'd1463;
            12'd366: current_page <= 12'd1985;
            12'd367: current_page <= 12'd454;
            12'd368: current_page <= 12'd976;
            12'd369: current_page <= 12'd1498;
            12'd370: current_page <= 12'd2020;
            12'd371: current_page <= 12'd489;
            12'd372: current_page <= 12'd1011;
            12'd373: current_page <= 12'd1533;
            12'd374: current_page <= 12'd2;
            12'd375: current_page <= 12'd524;
            12'd376: current_page <= 12'd1046;
            12'd377: current_page <= 12'd1568;
            12'd378: current_page <= 12'd37;
            12'd379: current_page <= 12'd559;
            12'd380: current_page <= 12'd1081;
            12'd381: current_page <= 12'd1603;
            12'd382: current_page <= 12'd72;
            12'd383: current_page <= 12'd594;
            12'd384: current_page <= 12'd1116;
            12'd385: current_page <= 12'd1638;
            12'd386: current_page <= 12'd107;
            12'd387: current_page <= 12'd629;
            12'd388: current_page <= 12'd1151;
            12'd389: current_page <= 12'd1673;
            12'd390: current_page <= 12'd142;
            12'd391: current_page <= 12'd664;
            12'd392: current_page <= 12'd1186;
            12'd393: current_page <= 12'd1708;
            12'd394: current_page <= 12'd177;
            12'd395: current_page <= 12'd699;
            12'd396: current_page <= 12'd1221;
            12'd397: current_page <= 12'd1743;
            12'd398: current_page <= 12'd212;
            12'd399: current_page <= 12'd734;
            12'd400: current_page <= 12'd1256;
            12'd401: current_page <= 12'd1778;
            12'd402: current_page <= 12'd247;
            12'd403: current_page <= 12'd769;
            12'd404: current_page <= 12'd1291;
            12'd405: current_page <= 12'd1813;
            12'd406: current_page <= 12'd282;
            12'd407: current_page <= 12'd804;
            12'd408: current_page <= 12'd1326;
            12'd409: current_page <= 12'd1848;
            12'd410: current_page <= 12'd317;
            12'd411: current_page <= 12'd839;
            12'd412: current_page <= 12'd1361;
            12'd413: current_page <= 12'd1883;
            12'd414: current_page <= 12'd352;
            12'd415: current_page <= 12'd874;
            12'd416: current_page <= 12'd1396;
            12'd417: current_page <= 12'd1918;
            12'd418: current_page <= 12'd387;
            12'd419: current_page <= 12'd909;
            12'd420: current_page <= 12'd1431;
            12'd421: current_page <= 12'd1953;
            12'd422: current_page <= 12'd422;
            12'd423: current_page <= 12'd944;
            12'd424: current_page <= 12'd1466;
            12'd425: current_page <= 12'd1988;
            12'd426: current_page <= 12'd457;
            12'd427: current_page <= 12'd979;
            12'd428: current_page <= 12'd1501;
            12'd429: current_page <= 12'd2023;
            12'd430: current_page <= 12'd492;
            12'd431: current_page <= 12'd1014;
            12'd432: current_page <= 12'd1536;
            12'd433: current_page <= 12'd5;
            12'd434: current_page <= 12'd527;
            12'd435: current_page <= 12'd1049;
            12'd436: current_page <= 12'd1571;
            12'd437: current_page <= 12'd40;
            12'd438: current_page <= 12'd562;
            12'd439: current_page <= 12'd1084;
            12'd440: current_page <= 12'd1606;
            12'd441: current_page <= 12'd75;
            12'd442: current_page <= 12'd597;
            12'd443: current_page <= 12'd1119;
            12'd444: current_page <= 12'd1641;
            12'd445: current_page <= 12'd110;
            12'd446: current_page <= 12'd632;
            12'd447: current_page <= 12'd1154;
            12'd448: current_page <= 12'd1676;
            12'd449: current_page <= 12'd145;
            12'd450: current_page <= 12'd667;
            12'd451: current_page <= 12'd1189;
            12'd452: current_page <= 12'd1711;
            12'd453: current_page <= 12'd180;
            12'd454: current_page <= 12'd702;
            12'd455: current_page <= 12'd1224;
            12'd456: current_page <= 12'd1746;
            12'd457: current_page <= 12'd215;
            12'd458: current_page <= 12'd737;
            12'd459: current_page <= 12'd1259;
            12'd460: current_page <= 12'd1781;
            12'd461: current_page <= 12'd250;
            12'd462: current_page <= 12'd772;
            12'd463: current_page <= 12'd1294;
            12'd464: current_page <= 12'd1816;
            12'd465: current_page <= 12'd285;
            12'd466: current_page <= 12'd807;
            12'd467: current_page <= 12'd1329;
            12'd468: current_page <= 12'd1851;
            12'd469: current_page <= 12'd320;
            12'd470: current_page <= 12'd842;
            12'd471: current_page <= 12'd1364;
            12'd472: current_page <= 12'd1886;
            12'd473: current_page <= 12'd355;
            12'd474: current_page <= 12'd877;
            12'd475: current_page <= 12'd1399;
            12'd476: current_page <= 12'd1921;
            12'd477: current_page <= 12'd390;
            12'd478: current_page <= 12'd912;
            12'd479: current_page <= 12'd1434;
            12'd480: current_page <= 12'd1956;
            12'd481: current_page <= 12'd425;
            12'd482: current_page <= 12'd947;
            12'd483: current_page <= 12'd1469;
            12'd484: current_page <= 12'd1991;
            12'd485: current_page <= 12'd460;
            12'd486: current_page <= 12'd982;
            12'd487: current_page <= 12'd1504;
            12'd488: current_page <= 12'd2026;
            12'd489: current_page <= 12'd495;
            12'd490: current_page <= 12'd1017;
            12'd491: current_page <= 12'd1539;
            12'd492: current_page <= 12'd8;
            12'd493: current_page <= 12'd530;
            12'd494: current_page <= 12'd1052;
            12'd495: current_page <= 12'd1574;
            12'd496: current_page <= 12'd43;
            12'd497: current_page <= 12'd565;
            12'd498: current_page <= 12'd1087;
            12'd499: current_page <= 12'd1609;
            12'd500: current_page <= 12'd78;
            12'd501: current_page <= 12'd600;
            12'd502: current_page <= 12'd1122;
            12'd503: current_page <= 12'd1644;
            12'd504: current_page <= 12'd113;
            12'd505: current_page <= 12'd635;
            12'd506: current_page <= 12'd1157;
            12'd507: current_page <= 12'd1679;
            12'd508: current_page <= 12'd148;
            12'd509: current_page <= 12'd670;
            12'd510: current_page <= 12'd1192;
            12'd511: current_page <= 12'd1714;
            12'd512: current_page <= 12'd183;
            12'd513: current_page <= 12'd705;
            12'd514: current_page <= 12'd1227;
            12'd515: current_page <= 12'd1749;
            12'd516: current_page <= 12'd218;
            12'd517: current_page <= 12'd740;
            12'd518: current_page <= 12'd1262;
            12'd519: current_page <= 12'd1784;
            12'd520: current_page <= 12'd253;
            12'd521: current_page <= 12'd775;
            12'd522: current_page <= 12'd1297;
            12'd523: current_page <= 12'd1819;
            12'd524: current_page <= 12'd288;
            12'd525: current_page <= 12'd810;
            12'd526: current_page <= 12'd1332;
            12'd527: current_page <= 12'd1854;
            12'd528: current_page <= 12'd323;
            12'd529: current_page <= 12'd845;
            12'd530: current_page <= 12'd1367;
            12'd531: current_page <= 12'd1889;
            12'd532: current_page <= 12'd358;
            12'd533: current_page <= 12'd880;
            12'd534: current_page <= 12'd1402;
            12'd535: current_page <= 12'd1924;
            12'd536: current_page <= 12'd393;
            12'd537: current_page <= 12'd915;
            12'd538: current_page <= 12'd1437;
            12'd539: current_page <= 12'd1959;
            12'd540: current_page <= 12'd428;
            12'd541: current_page <= 12'd950;
            12'd542: current_page <= 12'd1472;
            12'd543: current_page <= 12'd1994;
            12'd544: current_page <= 12'd463;
            12'd545: current_page <= 12'd985;
            12'd546: current_page <= 12'd1507;
            12'd547: current_page <= 12'd2029;
            12'd548: current_page <= 12'd498;
            12'd549: current_page <= 12'd1020;
            12'd550: current_page <= 12'd1542;
            12'd551: current_page <= 12'd11;
            12'd552: current_page <= 12'd533;
            12'd553: current_page <= 12'd1055;
            12'd554: current_page <= 12'd1577;
            12'd555: current_page <= 12'd46;
            12'd556: current_page <= 12'd568;
            12'd557: current_page <= 12'd1090;
            12'd558: current_page <= 12'd1612;
            12'd559: current_page <= 12'd81;
            12'd560: current_page <= 12'd603;
            12'd561: current_page <= 12'd1125;
            12'd562: current_page <= 12'd1647;
            12'd563: current_page <= 12'd116;
            12'd564: current_page <= 12'd638;
            12'd565: current_page <= 12'd1160;
            12'd566: current_page <= 12'd1682;
            12'd567: current_page <= 12'd151;
            12'd568: current_page <= 12'd673;
            12'd569: current_page <= 12'd1195;
            12'd570: current_page <= 12'd1717;
            12'd571: current_page <= 12'd186;
            12'd572: current_page <= 12'd708;
            12'd573: current_page <= 12'd1230;
            12'd574: current_page <= 12'd1752;
            12'd575: current_page <= 12'd221;
            12'd576: current_page <= 12'd743;
            12'd577: current_page <= 12'd1265;
            12'd578: current_page <= 12'd1787;
            12'd579: current_page <= 12'd256;
            12'd580: current_page <= 12'd778;
            12'd581: current_page <= 12'd1300;
            12'd582: current_page <= 12'd1822;
            12'd583: current_page <= 12'd291;
            12'd584: current_page <= 12'd813;
            12'd585: current_page <= 12'd1335;
            12'd586: current_page <= 12'd1857;
            12'd587: current_page <= 12'd326;
            12'd588: current_page <= 12'd848;
            12'd589: current_page <= 12'd1370;
            12'd590: current_page <= 12'd1892;
            12'd591: current_page <= 12'd361;
            12'd592: current_page <= 12'd883;
            12'd593: current_page <= 12'd1405;
            12'd594: current_page <= 12'd1927;
            12'd595: current_page <= 12'd396;
            12'd596: current_page <= 12'd918;
            12'd597: current_page <= 12'd1440;
            12'd598: current_page <= 12'd1962;
            12'd599: current_page <= 12'd431;
            12'd600: current_page <= 12'd953;
            12'd601: current_page <= 12'd1475;
            12'd602: current_page <= 12'd1997;
            12'd603: current_page <= 12'd466;
            12'd604: current_page <= 12'd988;
            12'd605: current_page <= 12'd1510;
            12'd606: current_page <= 12'd2032;
            12'd607: current_page <= 12'd501;
            12'd608: current_page <= 12'd1023;
            12'd609: current_page <= 12'd1545;
            12'd610: current_page <= 12'd14;
            12'd611: current_page <= 12'd536;
            12'd612: current_page <= 12'd1058;
            12'd613: current_page <= 12'd1580;
            12'd614: current_page <= 12'd49;
            12'd615: current_page <= 12'd571;
            12'd616: current_page <= 12'd1093;
            12'd617: current_page <= 12'd1615;
            12'd618: current_page <= 12'd84;
            12'd619: current_page <= 12'd606;
            12'd620: current_page <= 12'd1128;
            12'd621: current_page <= 12'd1650;
            12'd622: current_page <= 12'd119;
            12'd623: current_page <= 12'd641;
            12'd624: current_page <= 12'd1163;
            12'd625: current_page <= 12'd1685;
            12'd626: current_page <= 12'd154;
            12'd627: current_page <= 12'd676;
            12'd628: current_page <= 12'd1198;
            12'd629: current_page <= 12'd1720;
            12'd630: current_page <= 12'd189;
            12'd631: current_page <= 12'd711;
            12'd632: current_page <= 12'd1233;
            12'd633: current_page <= 12'd1755;
            12'd634: current_page <= 12'd224;
            12'd635: current_page <= 12'd746;
            12'd636: current_page <= 12'd1268;
            12'd637: current_page <= 12'd1790;
            12'd638: current_page <= 12'd259;
            12'd639: current_page <= 12'd781;
            12'd640: current_page <= 12'd1303;
            12'd641: current_page <= 12'd1825;
            12'd642: current_page <= 12'd294;
            12'd643: current_page <= 12'd816;
            12'd644: current_page <= 12'd1338;
            12'd645: current_page <= 12'd1860;
            12'd646: current_page <= 12'd329;
            12'd647: current_page <= 12'd851;
            12'd648: current_page <= 12'd1373;
            12'd649: current_page <= 12'd1895;
            12'd650: current_page <= 12'd364;
            12'd651: current_page <= 12'd886;
            12'd652: current_page <= 12'd1408;
            12'd653: current_page <= 12'd1930;
            12'd654: current_page <= 12'd399;
            12'd655: current_page <= 12'd921;
            12'd656: current_page <= 12'd1443;
            12'd657: current_page <= 12'd1965;
            12'd658: current_page <= 12'd434;
            12'd659: current_page <= 12'd956;
            12'd660: current_page <= 12'd1478;
            12'd661: current_page <= 12'd2000;
            12'd662: current_page <= 12'd469;
            12'd663: current_page <= 12'd991;
            12'd664: current_page <= 12'd1513;
            12'd665: current_page <= 12'd2035;
            12'd666: current_page <= 12'd504;
            12'd667: current_page <= 12'd1026;
            12'd668: current_page <= 12'd1548;
            12'd669: current_page <= 12'd17;
            12'd670: current_page <= 12'd539;
            12'd671: current_page <= 12'd1061;
            12'd672: current_page <= 12'd1583;
            12'd673: current_page <= 12'd52;
            12'd674: current_page <= 12'd574;
            12'd675: current_page <= 12'd1096;
            12'd676: current_page <= 12'd1618;
            12'd677: current_page <= 12'd87;
            12'd678: current_page <= 12'd609;
            12'd679: current_page <= 12'd1131;
            12'd680: current_page <= 12'd1653;
            12'd681: current_page <= 12'd122;
            12'd682: current_page <= 12'd644;
            12'd683: current_page <= 12'd1166;
            12'd684: current_page <= 12'd1688;
            12'd685: current_page <= 12'd157;
            12'd686: current_page <= 12'd679;
            12'd687: current_page <= 12'd1201;
            12'd688: current_page <= 12'd1723;
            12'd689: current_page <= 12'd192;
            12'd690: current_page <= 12'd714;
            12'd691: current_page <= 12'd1236;
            12'd692: current_page <= 12'd1758;
            12'd693: current_page <= 12'd227;
            12'd694: current_page <= 12'd749;
            12'd695: current_page <= 12'd1271;
            12'd696: current_page <= 12'd1793;
            12'd697: current_page <= 12'd262;
            12'd698: current_page <= 12'd784;
            12'd699: current_page <= 12'd1306;
            12'd700: current_page <= 12'd1828;
            12'd701: current_page <= 12'd297;
            12'd702: current_page <= 12'd819;
            12'd703: current_page <= 12'd1341;
            12'd704: current_page <= 12'd1863;
            12'd705: current_page <= 12'd332;
            12'd706: current_page <= 12'd854;
            12'd707: current_page <= 12'd1376;
            12'd708: current_page <= 12'd1898;
            12'd709: current_page <= 12'd367;
            12'd710: current_page <= 12'd889;
            12'd711: current_page <= 12'd1411;
            12'd712: current_page <= 12'd1933;
            12'd713: current_page <= 12'd402;
            12'd714: current_page <= 12'd924;
            12'd715: current_page <= 12'd1446;
            12'd716: current_page <= 12'd1968;
            12'd717: current_page <= 12'd437;
            12'd718: current_page <= 12'd959;
            12'd719: current_page <= 12'd1481;
            12'd720: current_page <= 12'd2003;
            12'd721: current_page <= 12'd472;
            12'd722: current_page <= 12'd994;
            12'd723: current_page <= 12'd1516;
            12'd724: current_page <= 12'd2038;
            12'd725: current_page <= 12'd507;
            12'd726: current_page <= 12'd1029;
            12'd727: current_page <= 12'd1551;
            12'd728: current_page <= 12'd20;
            12'd729: current_page <= 12'd542;
            12'd730: current_page <= 12'd1064;
            12'd731: current_page <= 12'd1586;
            12'd732: current_page <= 12'd55;
            12'd733: current_page <= 12'd577;
            12'd734: current_page <= 12'd1099;
            12'd735: current_page <= 12'd1621;
            12'd736: current_page <= 12'd90;
            12'd737: current_page <= 12'd612;
            12'd738: current_page <= 12'd1134;
            12'd739: current_page <= 12'd1656;
            12'd740: current_page <= 12'd125;
            12'd741: current_page <= 12'd647;
            12'd742: current_page <= 12'd1169;
            12'd743: current_page <= 12'd1691;
            12'd744: current_page <= 12'd160;
            12'd745: current_page <= 12'd682;
            12'd746: current_page <= 12'd1204;
            12'd747: current_page <= 12'd1726;
            12'd748: current_page <= 12'd195;
            12'd749: current_page <= 12'd717;
            12'd750: current_page <= 12'd1239;
            12'd751: current_page <= 12'd1761;
            12'd752: current_page <= 12'd230;
            12'd753: current_page <= 12'd752;
            12'd754: current_page <= 12'd1274;
            12'd755: current_page <= 12'd1796;
            12'd756: current_page <= 12'd265;
            12'd757: current_page <= 12'd787;
            12'd758: current_page <= 12'd1309;
            12'd759: current_page <= 12'd1831;
            12'd760: current_page <= 12'd300;
            12'd761: current_page <= 12'd822;
            12'd762: current_page <= 12'd1344;
            12'd763: current_page <= 12'd1866;
            12'd764: current_page <= 12'd335;
            12'd765: current_page <= 12'd857;
            12'd766: current_page <= 12'd1379;
            12'd767: current_page <= 12'd1901;
            12'd768: current_page <= 12'd370;
            12'd769: current_page <= 12'd892;
            12'd770: current_page <= 12'd1414;
            12'd771: current_page <= 12'd1936;
            12'd772: current_page <= 12'd405;
            12'd773: current_page <= 12'd927;
            12'd774: current_page <= 12'd1449;
            12'd775: current_page <= 12'd1971;
            12'd776: current_page <= 12'd440;
            12'd777: current_page <= 12'd962;
            12'd778: current_page <= 12'd1484;
            12'd779: current_page <= 12'd2006;
            12'd780: current_page <= 12'd475;
            12'd781: current_page <= 12'd997;
            12'd782: current_page <= 12'd1519;
            12'd783: current_page <= 12'd2041;
            12'd784: current_page <= 12'd510;
            12'd785: current_page <= 12'd1032;
            12'd786: current_page <= 12'd1554;
            12'd787: current_page <= 12'd23;
            12'd788: current_page <= 12'd545;
            12'd789: current_page <= 12'd1067;
            12'd790: current_page <= 12'd1589;
            12'd791: current_page <= 12'd58;
            12'd792: current_page <= 12'd580;
            12'd793: current_page <= 12'd1102;
            12'd794: current_page <= 12'd1624;
            12'd795: current_page <= 12'd93;
            12'd796: current_page <= 12'd615;
            12'd797: current_page <= 12'd1137;
            12'd798: current_page <= 12'd1659;
            12'd799: current_page <= 12'd128;
            12'd800: current_page <= 12'd650;
            12'd801: current_page <= 12'd1172;
            12'd802: current_page <= 12'd1694;
            12'd803: current_page <= 12'd163;
            12'd804: current_page <= 12'd685;
            12'd805: current_page <= 12'd1207;
            12'd806: current_page <= 12'd1729;
            12'd807: current_page <= 12'd198;
            12'd808: current_page <= 12'd720;
            12'd809: current_page <= 12'd1242;
            12'd810: current_page <= 12'd1764;
            12'd811: current_page <= 12'd233;
            12'd812: current_page <= 12'd755;
            12'd813: current_page <= 12'd1277;
            12'd814: current_page <= 12'd1799;
            12'd815: current_page <= 12'd268;
            12'd816: current_page <= 12'd790;
            12'd817: current_page <= 12'd1312;
            12'd818: current_page <= 12'd1834;
            12'd819: current_page <= 12'd303;
            12'd820: current_page <= 12'd825;
            12'd821: current_page <= 12'd1347;
            12'd822: current_page <= 12'd1869;
            12'd823: current_page <= 12'd338;
            12'd824: current_page <= 12'd860;
            12'd825: current_page <= 12'd1382;
            12'd826: current_page <= 12'd1904;
            12'd827: current_page <= 12'd373;
            12'd828: current_page <= 12'd895;
            12'd829: current_page <= 12'd1417;
            12'd830: current_page <= 12'd1939;
            12'd831: current_page <= 12'd408;
            12'd832: current_page <= 12'd930;
            12'd833: current_page <= 12'd1452;
            12'd834: current_page <= 12'd1974;
            12'd835: current_page <= 12'd443;
            12'd836: current_page <= 12'd965;
            12'd837: current_page <= 12'd1487;
            12'd838: current_page <= 12'd2009;
            12'd839: current_page <= 12'd478;
            12'd840: current_page <= 12'd1000;
            12'd841: current_page <= 12'd1522;
            12'd842: current_page <= 12'd2044;
            12'd843: current_page <= 12'd513;
            12'd844: current_page <= 12'd1035;
            12'd845: current_page <= 12'd1557;
            12'd846: current_page <= 12'd26;
            12'd847: current_page <= 12'd548;
            12'd848: current_page <= 12'd1070;
            12'd849: current_page <= 12'd1592;
            12'd850: current_page <= 12'd61;
            12'd851: current_page <= 12'd583;
            12'd852: current_page <= 12'd1105;
            12'd853: current_page <= 12'd1627;
            12'd854: current_page <= 12'd96;
            12'd855: current_page <= 12'd618;
            12'd856: current_page <= 12'd1140;
            12'd857: current_page <= 12'd1662;
            12'd858: current_page <= 12'd131;
            12'd859: current_page <= 12'd653;
            12'd860: current_page <= 12'd1175;
            12'd861: current_page <= 12'd1697;
            12'd862: current_page <= 12'd166;
            12'd863: current_page <= 12'd688;
            12'd864: current_page <= 12'd1210;
            12'd865: current_page <= 12'd1732;
            12'd866: current_page <= 12'd201;
            12'd867: current_page <= 12'd723;
            12'd868: current_page <= 12'd1245;
            12'd869: current_page <= 12'd1767;
            12'd870: current_page <= 12'd236;
            12'd871: current_page <= 12'd758;
            12'd872: current_page <= 12'd1280;
            12'd873: current_page <= 12'd1802;
            12'd874: current_page <= 12'd271;
            12'd875: current_page <= 12'd793;
            12'd876: current_page <= 12'd1315;
            12'd877: current_page <= 12'd1837;
            12'd878: current_page <= 12'd306;
            12'd879: current_page <= 12'd828;
            12'd880: current_page <= 12'd1350;
            12'd881: current_page <= 12'd1872;
            12'd882: current_page <= 12'd341;
            12'd883: current_page <= 12'd863;
            12'd884: current_page <= 12'd1385;
            12'd885: current_page <= 12'd1907;
            12'd886: current_page <= 12'd376;
            12'd887: current_page <= 12'd898;
            12'd888: current_page <= 12'd1420;
            12'd889: current_page <= 12'd1942;
            12'd890: current_page <= 12'd411;
            12'd891: current_page <= 12'd933;
            12'd892: current_page <= 12'd1455;
            12'd893: current_page <= 12'd1977;
            12'd894: current_page <= 12'd446;
            12'd895: current_page <= 12'd968;
            12'd896: current_page <= 12'd1490;
            12'd897: current_page <= 12'd2012;
            12'd898: current_page <= 12'd481;
            12'd899: current_page <= 12'd1003;
            12'd900: current_page <= 12'd1525;
            12'd901: current_page <= 12'd2047;
            12'd902: current_page <= 12'd516;
            12'd903: current_page <= 12'd1038;
            12'd904: current_page <= 12'd1560;
            12'd905: current_page <= 12'd29;
            12'd906: current_page <= 12'd551;
            12'd907: current_page <= 12'd1073;
            12'd908: current_page <= 12'd1595;
            12'd909: current_page <= 12'd64;
            12'd910: current_page <= 12'd586;
            12'd911: current_page <= 12'd1108;
            12'd912: current_page <= 12'd1630;
            12'd913: current_page <= 12'd99;
            12'd914: current_page <= 12'd621;
            12'd915: current_page <= 12'd1143;
            12'd916: current_page <= 12'd1665;
            12'd917: current_page <= 12'd134;
            12'd918: current_page <= 12'd656;
            12'd919: current_page <= 12'd1178;
            12'd920: current_page <= 12'd1700;
            12'd921: current_page <= 12'd169;
            12'd922: current_page <= 12'd691;
            12'd923: current_page <= 12'd1213;
            12'd924: current_page <= 12'd1735;
            12'd925: current_page <= 12'd204;
            12'd926: current_page <= 12'd726;
            12'd927: current_page <= 12'd1248;
            12'd928: current_page <= 12'd1770;
            12'd929: current_page <= 12'd239;
            12'd930: current_page <= 12'd761;
            12'd931: current_page <= 12'd1283;
            12'd932: current_page <= 12'd1805;
            12'd933: current_page <= 12'd274;
            12'd934: current_page <= 12'd796;
            12'd935: current_page <= 12'd1318;
            12'd936: current_page <= 12'd1840;
            12'd937: current_page <= 12'd309;
            12'd938: current_page <= 12'd831;
            12'd939: current_page <= 12'd1353;
            12'd940: current_page <= 12'd1875;
            12'd941: current_page <= 12'd344;
            12'd942: current_page <= 12'd866;
            12'd943: current_page <= 12'd1388;
            12'd944: current_page <= 12'd1910;
            12'd945: current_page <= 12'd379;
            12'd946: current_page <= 12'd901;
            12'd947: current_page <= 12'd1423;
            12'd948: current_page <= 12'd1945;
            12'd949: current_page <= 12'd414;
            12'd950: current_page <= 12'd936;
            12'd951: current_page <= 12'd1458;
            12'd952: current_page <= 12'd1980;
            12'd953: current_page <= 12'd449;
            12'd954: current_page <= 12'd971;
            12'd955: current_page <= 12'd1493;
            12'd956: current_page <= 12'd2015;
            12'd957: current_page <= 12'd484;
            12'd958: current_page <= 12'd1006;
            12'd959: current_page <= 12'd1528;
            12'd960: current_page <= 12'd2050;
            12'd961: current_page <= 12'd519;
            12'd962: current_page <= 12'd1041;
            12'd963: current_page <= 12'd1563;
            12'd964: current_page <= 12'd32;
            12'd965: current_page <= 12'd554;
            12'd966: current_page <= 12'd1076;
            12'd967: current_page <= 12'd1598;
            12'd968: current_page <= 12'd67;
            12'd969: current_page <= 12'd589;
            12'd970: current_page <= 12'd1111;
            12'd971: current_page <= 12'd1633;
            12'd972: current_page <= 12'd102;
            12'd973: current_page <= 12'd624;
            12'd974: current_page <= 12'd1146;
            12'd975: current_page <= 12'd1668;
            12'd976: current_page <= 12'd137;
            12'd977: current_page <= 12'd659;
            12'd978: current_page <= 12'd1181;
            12'd979: current_page <= 12'd1703;
            12'd980: current_page <= 12'd172;
            12'd981: current_page <= 12'd694;
            12'd982: current_page <= 12'd1216;
            12'd983: current_page <= 12'd1738;
            12'd984: current_page <= 12'd207;
            12'd985: current_page <= 12'd729;
            12'd986: current_page <= 12'd1251;
            12'd987: current_page <= 12'd1773;
            12'd988: current_page <= 12'd242;
            12'd989: current_page <= 12'd764;
            12'd990: current_page <= 12'd1286;
            12'd991: current_page <= 12'd1808;
            12'd992: current_page <= 12'd277;
            12'd993: current_page <= 12'd799;
            12'd994: current_page <= 12'd1321;
            12'd995: current_page <= 12'd1843;
            12'd996: current_page <= 12'd312;
            12'd997: current_page <= 12'd834;
            12'd998: current_page <= 12'd1356;
            12'd999: current_page <= 12'd1878;
            12'd1000: current_page <= 12'd347;
            12'd1001: current_page <= 12'd869;
            12'd1002: current_page <= 12'd1391;
            12'd1003: current_page <= 12'd1913;
            12'd1004: current_page <= 12'd382;
            12'd1005: current_page <= 12'd904;
            12'd1006: current_page <= 12'd1426;
            12'd1007: current_page <= 12'd1948;
            12'd1008: current_page <= 12'd417;
            12'd1009: current_page <= 12'd939;
            12'd1010: current_page <= 12'd1461;
            12'd1011: current_page <= 12'd1983;
            12'd1012: current_page <= 12'd452;
            12'd1013: current_page <= 12'd974;
            12'd1014: current_page <= 12'd1496;
            12'd1015: current_page <= 12'd2018;
            12'd1016: current_page <= 12'd487;
            12'd1017: current_page <= 12'd1009;
            12'd1018: current_page <= 12'd1531;
            12'd1019: current_page <= 12'd0;
            12'd1020: current_page <= 12'd522;
            12'd1021: current_page <= 12'd1044;
            12'd1022: current_page <= 12'd1566;
            12'd1023: current_page <= 12'd35;
            12'd1024: current_page <= 12'd557;
            12'd1025: current_page <= 12'd1079;
            12'd1026: current_page <= 12'd1601;
            12'd1027: current_page <= 12'd70;
            12'd1028: current_page <= 12'd592;
            12'd1029: current_page <= 12'd1114;
            12'd1030: current_page <= 12'd1636;
            12'd1031: current_page <= 12'd105;
            12'd1032: current_page <= 12'd627;
            12'd1033: current_page <= 12'd1149;
            12'd1034: current_page <= 12'd1671;
            12'd1035: current_page <= 12'd140;
            12'd1036: current_page <= 12'd662;
            12'd1037: current_page <= 12'd1184;
            12'd1038: current_page <= 12'd1706;
            12'd1039: current_page <= 12'd175;
            12'd1040: current_page <= 12'd697;
            12'd1041: current_page <= 12'd1219;
            12'd1042: current_page <= 12'd1741;
            12'd1043: current_page <= 12'd210;
            12'd1044: current_page <= 12'd732;
            12'd1045: current_page <= 12'd1254;
            12'd1046: current_page <= 12'd1776;
            12'd1047: current_page <= 12'd245;
            12'd1048: current_page <= 12'd767;
            12'd1049: current_page <= 12'd1289;
            12'd1050: current_page <= 12'd1811;
            12'd1051: current_page <= 12'd280;
            12'd1052: current_page <= 12'd802;
            12'd1053: current_page <= 12'd1324;
            12'd1054: current_page <= 12'd1846;
            12'd1055: current_page <= 12'd315;
            12'd1056: current_page <= 12'd837;
            12'd1057: current_page <= 12'd1359;
            12'd1058: current_page <= 12'd1881;
            12'd1059: current_page <= 12'd350;
            12'd1060: current_page <= 12'd872;
            12'd1061: current_page <= 12'd1394;
            12'd1062: current_page <= 12'd1916;
            12'd1063: current_page <= 12'd385;
            12'd1064: current_page <= 12'd907;
            12'd1065: current_page <= 12'd1429;
            12'd1066: current_page <= 12'd1951;
            12'd1067: current_page <= 12'd420;
            12'd1068: current_page <= 12'd942;
            12'd1069: current_page <= 12'd1464;
            12'd1070: current_page <= 12'd1986;
            12'd1071: current_page <= 12'd455;
            12'd1072: current_page <= 12'd977;
            12'd1073: current_page <= 12'd1499;
            12'd1074: current_page <= 12'd2021;
            12'd1075: current_page <= 12'd490;
            12'd1076: current_page <= 12'd1012;
            12'd1077: current_page <= 12'd1534;
            12'd1078: current_page <= 12'd3;
            12'd1079: current_page <= 12'd525;
            12'd1080: current_page <= 12'd1047;
            12'd1081: current_page <= 12'd1569;
            12'd1082: current_page <= 12'd38;
            12'd1083: current_page <= 12'd560;
            12'd1084: current_page <= 12'd1082;
            12'd1085: current_page <= 12'd1604;
            12'd1086: current_page <= 12'd73;
            12'd1087: current_page <= 12'd595;
            12'd1088: current_page <= 12'd1117;
            12'd1089: current_page <= 12'd1639;
            12'd1090: current_page <= 12'd108;
            12'd1091: current_page <= 12'd630;
            12'd1092: current_page <= 12'd1152;
            12'd1093: current_page <= 12'd1674;
            12'd1094: current_page <= 12'd143;
            12'd1095: current_page <= 12'd665;
            12'd1096: current_page <= 12'd1187;
            12'd1097: current_page <= 12'd1709;
            12'd1098: current_page <= 12'd178;
            12'd1099: current_page <= 12'd700;
            12'd1100: current_page <= 12'd1222;
            12'd1101: current_page <= 12'd1744;
            12'd1102: current_page <= 12'd213;
            12'd1103: current_page <= 12'd735;
            12'd1104: current_page <= 12'd1257;
            12'd1105: current_page <= 12'd1779;
            12'd1106: current_page <= 12'd248;
            12'd1107: current_page <= 12'd770;
            12'd1108: current_page <= 12'd1292;
            12'd1109: current_page <= 12'd1814;
            12'd1110: current_page <= 12'd283;
            12'd1111: current_page <= 12'd805;
            12'd1112: current_page <= 12'd1327;
            12'd1113: current_page <= 12'd1849;
            12'd1114: current_page <= 12'd318;
            12'd1115: current_page <= 12'd840;
            12'd1116: current_page <= 12'd1362;
            12'd1117: current_page <= 12'd1884;
            12'd1118: current_page <= 12'd353;
            12'd1119: current_page <= 12'd875;
            12'd1120: current_page <= 12'd1397;
            12'd1121: current_page <= 12'd1919;
            12'd1122: current_page <= 12'd388;
            12'd1123: current_page <= 12'd910;
            12'd1124: current_page <= 12'd1432;
            12'd1125: current_page <= 12'd1954;
            12'd1126: current_page <= 12'd423;
            12'd1127: current_page <= 12'd945;
            12'd1128: current_page <= 12'd1467;
            12'd1129: current_page <= 12'd1989;
            12'd1130: current_page <= 12'd458;
            12'd1131: current_page <= 12'd980;
            12'd1132: current_page <= 12'd1502;
            12'd1133: current_page <= 12'd2024;
            12'd1134: current_page <= 12'd493;
            12'd1135: current_page <= 12'd1015;
            12'd1136: current_page <= 12'd1537;
            12'd1137: current_page <= 12'd6;
            12'd1138: current_page <= 12'd528;
            12'd1139: current_page <= 12'd1050;
            12'd1140: current_page <= 12'd1572;
            12'd1141: current_page <= 12'd41;
            12'd1142: current_page <= 12'd563;
            12'd1143: current_page <= 12'd1085;
            12'd1144: current_page <= 12'd1607;
            12'd1145: current_page <= 12'd76;
            12'd1146: current_page <= 12'd598;
            12'd1147: current_page <= 12'd1120;
            12'd1148: current_page <= 12'd1642;
            12'd1149: current_page <= 12'd111;
            12'd1150: current_page <= 12'd633;
            12'd1151: current_page <= 12'd1155;
            12'd1152: current_page <= 12'd1677;
            12'd1153: current_page <= 12'd146;
            12'd1154: current_page <= 12'd668;
            12'd1155: current_page <= 12'd1190;
            12'd1156: current_page <= 12'd1712;
            12'd1157: current_page <= 12'd181;
            12'd1158: current_page <= 12'd703;
            12'd1159: current_page <= 12'd1225;
            12'd1160: current_page <= 12'd1747;
            12'd1161: current_page <= 12'd216;
            12'd1162: current_page <= 12'd738;
            12'd1163: current_page <= 12'd1260;
            12'd1164: current_page <= 12'd1782;
            12'd1165: current_page <= 12'd251;
            12'd1166: current_page <= 12'd773;
            12'd1167: current_page <= 12'd1295;
            12'd1168: current_page <= 12'd1817;
            12'd1169: current_page <= 12'd286;
            12'd1170: current_page <= 12'd808;
            12'd1171: current_page <= 12'd1330;
            12'd1172: current_page <= 12'd1852;
            12'd1173: current_page <= 12'd321;
            12'd1174: current_page <= 12'd843;
            12'd1175: current_page <= 12'd1365;
            12'd1176: current_page <= 12'd1887;
            12'd1177: current_page <= 12'd356;
            12'd1178: current_page <= 12'd878;
            12'd1179: current_page <= 12'd1400;
            12'd1180: current_page <= 12'd1922;
            12'd1181: current_page <= 12'd391;
            12'd1182: current_page <= 12'd913;
            12'd1183: current_page <= 12'd1435;
            12'd1184: current_page <= 12'd1957;
            12'd1185: current_page <= 12'd426;
            12'd1186: current_page <= 12'd948;
            12'd1187: current_page <= 12'd1470;
            12'd1188: current_page <= 12'd1992;
            12'd1189: current_page <= 12'd461;
            12'd1190: current_page <= 12'd983;
            12'd1191: current_page <= 12'd1505;
            12'd1192: current_page <= 12'd2027;
            12'd1193: current_page <= 12'd496;
            12'd1194: current_page <= 12'd1018;
            12'd1195: current_page <= 12'd1540;
            12'd1196: current_page <= 12'd9;
            12'd1197: current_page <= 12'd531;
            12'd1198: current_page <= 12'd1053;
            12'd1199: current_page <= 12'd1575;
            12'd1200: current_page <= 12'd44;
            12'd1201: current_page <= 12'd566;
            12'd1202: current_page <= 12'd1088;
            12'd1203: current_page <= 12'd1610;
            12'd1204: current_page <= 12'd79;
            12'd1205: current_page <= 12'd601;
            12'd1206: current_page <= 12'd1123;
            12'd1207: current_page <= 12'd1645;
            12'd1208: current_page <= 12'd114;
            12'd1209: current_page <= 12'd636;
            12'd1210: current_page <= 12'd1158;
            12'd1211: current_page <= 12'd1680;
            12'd1212: current_page <= 12'd149;
            12'd1213: current_page <= 12'd671;
            12'd1214: current_page <= 12'd1193;
            12'd1215: current_page <= 12'd1715;
            12'd1216: current_page <= 12'd184;
            12'd1217: current_page <= 12'd706;
            12'd1218: current_page <= 12'd1228;
            12'd1219: current_page <= 12'd1750;
            12'd1220: current_page <= 12'd219;
            12'd1221: current_page <= 12'd741;
            12'd1222: current_page <= 12'd1263;
            12'd1223: current_page <= 12'd1785;
            12'd1224: current_page <= 12'd254;
            12'd1225: current_page <= 12'd776;
            12'd1226: current_page <= 12'd1298;
            12'd1227: current_page <= 12'd1820;
            12'd1228: current_page <= 12'd289;
            12'd1229: current_page <= 12'd811;
            12'd1230: current_page <= 12'd1333;
            12'd1231: current_page <= 12'd1855;
            12'd1232: current_page <= 12'd324;
            12'd1233: current_page <= 12'd846;
            12'd1234: current_page <= 12'd1368;
            12'd1235: current_page <= 12'd1890;
            12'd1236: current_page <= 12'd359;
            12'd1237: current_page <= 12'd881;
            12'd1238: current_page <= 12'd1403;
            12'd1239: current_page <= 12'd1925;
            12'd1240: current_page <= 12'd394;
            12'd1241: current_page <= 12'd916;
            12'd1242: current_page <= 12'd1438;
            12'd1243: current_page <= 12'd1960;
            12'd1244: current_page <= 12'd429;
            12'd1245: current_page <= 12'd951;
            12'd1246: current_page <= 12'd1473;
            12'd1247: current_page <= 12'd1995;
            12'd1248: current_page <= 12'd464;
            12'd1249: current_page <= 12'd986;
            12'd1250: current_page <= 12'd1508;
            12'd1251: current_page <= 12'd2030;
            12'd1252: current_page <= 12'd499;
            12'd1253: current_page <= 12'd1021;
            12'd1254: current_page <= 12'd1543;
            12'd1255: current_page <= 12'd12;
            12'd1256: current_page <= 12'd534;
            12'd1257: current_page <= 12'd1056;
            12'd1258: current_page <= 12'd1578;
            12'd1259: current_page <= 12'd47;
            12'd1260: current_page <= 12'd569;
            12'd1261: current_page <= 12'd1091;
            12'd1262: current_page <= 12'd1613;
            12'd1263: current_page <= 12'd82;
            12'd1264: current_page <= 12'd604;
            12'd1265: current_page <= 12'd1126;
            12'd1266: current_page <= 12'd1648;
            12'd1267: current_page <= 12'd117;
            12'd1268: current_page <= 12'd639;
            12'd1269: current_page <= 12'd1161;
            12'd1270: current_page <= 12'd1683;
            12'd1271: current_page <= 12'd152;
            12'd1272: current_page <= 12'd674;
            12'd1273: current_page <= 12'd1196;
            12'd1274: current_page <= 12'd1718;
            12'd1275: current_page <= 12'd187;
            12'd1276: current_page <= 12'd709;
            12'd1277: current_page <= 12'd1231;
            12'd1278: current_page <= 12'd1753;
            12'd1279: current_page <= 12'd222;
            12'd1280: current_page <= 12'd744;
            12'd1281: current_page <= 12'd1266;
            12'd1282: current_page <= 12'd1788;
            12'd1283: current_page <= 12'd257;
            12'd1284: current_page <= 12'd779;
            12'd1285: current_page <= 12'd1301;
            12'd1286: current_page <= 12'd1823;
            12'd1287: current_page <= 12'd292;
            12'd1288: current_page <= 12'd814;
            12'd1289: current_page <= 12'd1336;
            12'd1290: current_page <= 12'd1858;
            12'd1291: current_page <= 12'd327;
            12'd1292: current_page <= 12'd849;
            12'd1293: current_page <= 12'd1371;
            12'd1294: current_page <= 12'd1893;
            12'd1295: current_page <= 12'd362;
            12'd1296: current_page <= 12'd884;
            12'd1297: current_page <= 12'd1406;
            12'd1298: current_page <= 12'd1928;
            12'd1299: current_page <= 12'd397;
            12'd1300: current_page <= 12'd919;
            12'd1301: current_page <= 12'd1441;
            12'd1302: current_page <= 12'd1963;
            12'd1303: current_page <= 12'd432;
            12'd1304: current_page <= 12'd954;
            12'd1305: current_page <= 12'd1476;
            12'd1306: current_page <= 12'd1998;
            12'd1307: current_page <= 12'd467;
            12'd1308: current_page <= 12'd989;
            12'd1309: current_page <= 12'd1511;
            12'd1310: current_page <= 12'd2033;
            12'd1311: current_page <= 12'd502;
            12'd1312: current_page <= 12'd1024;
            12'd1313: current_page <= 12'd1546;
            12'd1314: current_page <= 12'd15;
            12'd1315: current_page <= 12'd537;
            12'd1316: current_page <= 12'd1059;
            12'd1317: current_page <= 12'd1581;
            12'd1318: current_page <= 12'd50;
            12'd1319: current_page <= 12'd572;
            12'd1320: current_page <= 12'd1094;
            12'd1321: current_page <= 12'd1616;
            12'd1322: current_page <= 12'd85;
            12'd1323: current_page <= 12'd607;
            12'd1324: current_page <= 12'd1129;
            12'd1325: current_page <= 12'd1651;
            12'd1326: current_page <= 12'd120;
            12'd1327: current_page <= 12'd642;
            12'd1328: current_page <= 12'd1164;
            12'd1329: current_page <= 12'd1686;
            12'd1330: current_page <= 12'd155;
            12'd1331: current_page <= 12'd677;
            12'd1332: current_page <= 12'd1199;
            12'd1333: current_page <= 12'd1721;
            12'd1334: current_page <= 12'd190;
            12'd1335: current_page <= 12'd712;
            12'd1336: current_page <= 12'd1234;
            12'd1337: current_page <= 12'd1756;
            12'd1338: current_page <= 12'd225;
            12'd1339: current_page <= 12'd747;
            12'd1340: current_page <= 12'd1269;
            12'd1341: current_page <= 12'd1791;
            12'd1342: current_page <= 12'd260;
            12'd1343: current_page <= 12'd782;
            12'd1344: current_page <= 12'd1304;
            12'd1345: current_page <= 12'd1826;
            12'd1346: current_page <= 12'd295;
            12'd1347: current_page <= 12'd817;
            12'd1348: current_page <= 12'd1339;
            12'd1349: current_page <= 12'd1861;
            12'd1350: current_page <= 12'd330;
            12'd1351: current_page <= 12'd852;
            12'd1352: current_page <= 12'd1374;
            12'd1353: current_page <= 12'd1896;
            12'd1354: current_page <= 12'd365;
            12'd1355: current_page <= 12'd887;
            12'd1356: current_page <= 12'd1409;
            12'd1357: current_page <= 12'd1931;
            12'd1358: current_page <= 12'd400;
            12'd1359: current_page <= 12'd922;
            12'd1360: current_page <= 12'd1444;
            12'd1361: current_page <= 12'd1966;
            12'd1362: current_page <= 12'd435;
            12'd1363: current_page <= 12'd957;
            12'd1364: current_page <= 12'd1479;
            12'd1365: current_page <= 12'd2001;
            12'd1366: current_page <= 12'd470;
            12'd1367: current_page <= 12'd992;
            12'd1368: current_page <= 12'd1514;
            12'd1369: current_page <= 12'd2036;
            12'd1370: current_page <= 12'd505;
            12'd1371: current_page <= 12'd1027;
            12'd1372: current_page <= 12'd1549;
            12'd1373: current_page <= 12'd18;
            12'd1374: current_page <= 12'd540;
            12'd1375: current_page <= 12'd1062;
            12'd1376: current_page <= 12'd1584;
            12'd1377: current_page <= 12'd53;
            12'd1378: current_page <= 12'd575;
            12'd1379: current_page <= 12'd1097;
            12'd1380: current_page <= 12'd1619;
            12'd1381: current_page <= 12'd88;
            12'd1382: current_page <= 12'd610;
            12'd1383: current_page <= 12'd1132;
            12'd1384: current_page <= 12'd1654;
            12'd1385: current_page <= 12'd123;
            12'd1386: current_page <= 12'd645;
            12'd1387: current_page <= 12'd1167;
            12'd1388: current_page <= 12'd1689;
            12'd1389: current_page <= 12'd158;
            12'd1390: current_page <= 12'd680;
            12'd1391: current_page <= 12'd1202;
            12'd1392: current_page <= 12'd1724;
            12'd1393: current_page <= 12'd193;
            12'd1394: current_page <= 12'd715;
            12'd1395: current_page <= 12'd1237;
            12'd1396: current_page <= 12'd1759;
            12'd1397: current_page <= 12'd228;
            12'd1398: current_page <= 12'd750;
            12'd1399: current_page <= 12'd1272;
            12'd1400: current_page <= 12'd1794;
            12'd1401: current_page <= 12'd263;
            12'd1402: current_page <= 12'd785;
            12'd1403: current_page <= 12'd1307;
            12'd1404: current_page <= 12'd1829;
            12'd1405: current_page <= 12'd298;
            12'd1406: current_page <= 12'd820;
            12'd1407: current_page <= 12'd1342;
            12'd1408: current_page <= 12'd1864;
            12'd1409: current_page <= 12'd333;
            12'd1410: current_page <= 12'd855;
            12'd1411: current_page <= 12'd1377;
            12'd1412: current_page <= 12'd1899;
            12'd1413: current_page <= 12'd368;
            12'd1414: current_page <= 12'd890;
            12'd1415: current_page <= 12'd1412;
            12'd1416: current_page <= 12'd1934;
            12'd1417: current_page <= 12'd403;
            12'd1418: current_page <= 12'd925;
            12'd1419: current_page <= 12'd1447;
            12'd1420: current_page <= 12'd1969;
            12'd1421: current_page <= 12'd438;
            12'd1422: current_page <= 12'd960;
            12'd1423: current_page <= 12'd1482;
            12'd1424: current_page <= 12'd2004;
            12'd1425: current_page <= 12'd473;
            12'd1426: current_page <= 12'd995;
            12'd1427: current_page <= 12'd1517;
            12'd1428: current_page <= 12'd2039;
            12'd1429: current_page <= 12'd508;
            12'd1430: current_page <= 12'd1030;
            12'd1431: current_page <= 12'd1552;
            12'd1432: current_page <= 12'd21;
            12'd1433: current_page <= 12'd543;
            12'd1434: current_page <= 12'd1065;
            12'd1435: current_page <= 12'd1587;
            12'd1436: current_page <= 12'd56;
            12'd1437: current_page <= 12'd578;
            12'd1438: current_page <= 12'd1100;
            12'd1439: current_page <= 12'd1622;
            12'd1440: current_page <= 12'd91;
            12'd1441: current_page <= 12'd613;
            12'd1442: current_page <= 12'd1135;
            12'd1443: current_page <= 12'd1657;
            12'd1444: current_page <= 12'd126;
            12'd1445: current_page <= 12'd648;
            12'd1446: current_page <= 12'd1170;
            12'd1447: current_page <= 12'd1692;
            12'd1448: current_page <= 12'd161;
            12'd1449: current_page <= 12'd683;
            12'd1450: current_page <= 12'd1205;
            12'd1451: current_page <= 12'd1727;
            12'd1452: current_page <= 12'd196;
            12'd1453: current_page <= 12'd718;
            12'd1454: current_page <= 12'd1240;
            12'd1455: current_page <= 12'd1762;
            12'd1456: current_page <= 12'd231;
            12'd1457: current_page <= 12'd753;
            12'd1458: current_page <= 12'd1275;
            12'd1459: current_page <= 12'd1797;
            12'd1460: current_page <= 12'd266;
            12'd1461: current_page <= 12'd788;
            12'd1462: current_page <= 12'd1310;
            12'd1463: current_page <= 12'd1832;
            12'd1464: current_page <= 12'd301;
            12'd1465: current_page <= 12'd823;
            12'd1466: current_page <= 12'd1345;
            12'd1467: current_page <= 12'd1867;
            12'd1468: current_page <= 12'd336;
            12'd1469: current_page <= 12'd858;
            12'd1470: current_page <= 12'd1380;
            12'd1471: current_page <= 12'd1902;
            12'd1472: current_page <= 12'd371;
            12'd1473: current_page <= 12'd893;
            12'd1474: current_page <= 12'd1415;
            12'd1475: current_page <= 12'd1937;
            12'd1476: current_page <= 12'd406;
            12'd1477: current_page <= 12'd928;
            12'd1478: current_page <= 12'd1450;
            12'd1479: current_page <= 12'd1972;
            12'd1480: current_page <= 12'd441;
            12'd1481: current_page <= 12'd963;
            12'd1482: current_page <= 12'd1485;
            12'd1483: current_page <= 12'd2007;
            12'd1484: current_page <= 12'd476;
            12'd1485: current_page <= 12'd998;
            12'd1486: current_page <= 12'd1520;
            12'd1487: current_page <= 12'd2042;
            12'd1488: current_page <= 12'd511;
            12'd1489: current_page <= 12'd1033;
            12'd1490: current_page <= 12'd1555;
            12'd1491: current_page <= 12'd24;
            12'd1492: current_page <= 12'd546;
            12'd1493: current_page <= 12'd1068;
            12'd1494: current_page <= 12'd1590;
            12'd1495: current_page <= 12'd59;
            12'd1496: current_page <= 12'd581;
            12'd1497: current_page <= 12'd1103;
            12'd1498: current_page <= 12'd1625;
            12'd1499: current_page <= 12'd94;
            12'd1500: current_page <= 12'd616;
            12'd1501: current_page <= 12'd1138;
            12'd1502: current_page <= 12'd1660;
            12'd1503: current_page <= 12'd129;
            12'd1504: current_page <= 12'd651;
            12'd1505: current_page <= 12'd1173;
            12'd1506: current_page <= 12'd1695;
            12'd1507: current_page <= 12'd164;
            12'd1508: current_page <= 12'd686;
            12'd1509: current_page <= 12'd1208;
            12'd1510: current_page <= 12'd1730;
            12'd1511: current_page <= 12'd199;
            12'd1512: current_page <= 12'd721;
            12'd1513: current_page <= 12'd1243;
            12'd1514: current_page <= 12'd1765;
            12'd1515: current_page <= 12'd234;
            12'd1516: current_page <= 12'd756;
            12'd1517: current_page <= 12'd1278;
            12'd1518: current_page <= 12'd1800;
            12'd1519: current_page <= 12'd269;
            12'd1520: current_page <= 12'd791;
            12'd1521: current_page <= 12'd1313;
            12'd1522: current_page <= 12'd1835;
            12'd1523: current_page <= 12'd304;
            12'd1524: current_page <= 12'd826;
            12'd1525: current_page <= 12'd1348;
            12'd1526: current_page <= 12'd1870;
            12'd1527: current_page <= 12'd339;
            12'd1528: current_page <= 12'd861;
            12'd1529: current_page <= 12'd1383;
            12'd1530: current_page <= 12'd1905;
            12'd1531: current_page <= 12'd374;
            12'd1532: current_page <= 12'd896;
            12'd1533: current_page <= 12'd1418;
            12'd1534: current_page <= 12'd1940;
            12'd1535: current_page <= 12'd409;
            12'd1536: current_page <= 12'd931;
            12'd1537: current_page <= 12'd1453;
            12'd1538: current_page <= 12'd1975;
            12'd1539: current_page <= 12'd444;
            12'd1540: current_page <= 12'd966;
            12'd1541: current_page <= 12'd1488;
            12'd1542: current_page <= 12'd2010;
            12'd1543: current_page <= 12'd479;
            12'd1544: current_page <= 12'd1001;
            12'd1545: current_page <= 12'd1523;
            12'd1546: current_page <= 12'd2045;
            12'd1547: current_page <= 12'd514;
            12'd1548: current_page <= 12'd1036;
            12'd1549: current_page <= 12'd1558;
            12'd1550: current_page <= 12'd27;
            12'd1551: current_page <= 12'd549;
            12'd1552: current_page <= 12'd1071;
            12'd1553: current_page <= 12'd1593;
            12'd1554: current_page <= 12'd62;
            12'd1555: current_page <= 12'd584;
            12'd1556: current_page <= 12'd1106;
            12'd1557: current_page <= 12'd1628;
            12'd1558: current_page <= 12'd97;
            12'd1559: current_page <= 12'd619;
            12'd1560: current_page <= 12'd1141;
            12'd1561: current_page <= 12'd1663;
            12'd1562: current_page <= 12'd132;
            12'd1563: current_page <= 12'd654;
            12'd1564: current_page <= 12'd1176;
            12'd1565: current_page <= 12'd1698;
            12'd1566: current_page <= 12'd167;
            12'd1567: current_page <= 12'd689;
            12'd1568: current_page <= 12'd1211;
            12'd1569: current_page <= 12'd1733;
            12'd1570: current_page <= 12'd202;
            12'd1571: current_page <= 12'd724;
            12'd1572: current_page <= 12'd1246;
            12'd1573: current_page <= 12'd1768;
            12'd1574: current_page <= 12'd237;
            12'd1575: current_page <= 12'd759;
            12'd1576: current_page <= 12'd1281;
            12'd1577: current_page <= 12'd1803;
            12'd1578: current_page <= 12'd272;
            12'd1579: current_page <= 12'd794;
            12'd1580: current_page <= 12'd1316;
            12'd1581: current_page <= 12'd1838;
            12'd1582: current_page <= 12'd307;
            12'd1583: current_page <= 12'd829;
            12'd1584: current_page <= 12'd1351;
            12'd1585: current_page <= 12'd1873;
            12'd1586: current_page <= 12'd342;
            12'd1587: current_page <= 12'd864;
            12'd1588: current_page <= 12'd1386;
            12'd1589: current_page <= 12'd1908;
            12'd1590: current_page <= 12'd377;
            12'd1591: current_page <= 12'd899;
            12'd1592: current_page <= 12'd1421;
            12'd1593: current_page <= 12'd1943;
            12'd1594: current_page <= 12'd412;
            12'd1595: current_page <= 12'd934;
            12'd1596: current_page <= 12'd1456;
            12'd1597: current_page <= 12'd1978;
            12'd1598: current_page <= 12'd447;
            12'd1599: current_page <= 12'd969;
            12'd1600: current_page <= 12'd1491;
            12'd1601: current_page <= 12'd2013;
            12'd1602: current_page <= 12'd482;
            12'd1603: current_page <= 12'd1004;
            12'd1604: current_page <= 12'd1526;
            12'd1605: current_page <= 12'd2048;
            12'd1606: current_page <= 12'd517;
            12'd1607: current_page <= 12'd1039;
            12'd1608: current_page <= 12'd1561;
            12'd1609: current_page <= 12'd30;
            12'd1610: current_page <= 12'd552;
            12'd1611: current_page <= 12'd1074;
            12'd1612: current_page <= 12'd1596;
            12'd1613: current_page <= 12'd65;
            12'd1614: current_page <= 12'd587;
            12'd1615: current_page <= 12'd1109;
            12'd1616: current_page <= 12'd1631;
            12'd1617: current_page <= 12'd100;
            12'd1618: current_page <= 12'd622;
            12'd1619: current_page <= 12'd1144;
            12'd1620: current_page <= 12'd1666;
            12'd1621: current_page <= 12'd135;
            12'd1622: current_page <= 12'd657;
            12'd1623: current_page <= 12'd1179;
            12'd1624: current_page <= 12'd1701;
            12'd1625: current_page <= 12'd170;
            12'd1626: current_page <= 12'd692;
            12'd1627: current_page <= 12'd1214;
            12'd1628: current_page <= 12'd1736;
            12'd1629: current_page <= 12'd205;
            12'd1630: current_page <= 12'd727;
            12'd1631: current_page <= 12'd1249;
            12'd1632: current_page <= 12'd1771;
            12'd1633: current_page <= 12'd240;
            12'd1634: current_page <= 12'd762;
            12'd1635: current_page <= 12'd1284;
            12'd1636: current_page <= 12'd1806;
            12'd1637: current_page <= 12'd275;
            12'd1638: current_page <= 12'd797;
            12'd1639: current_page <= 12'd1319;
            12'd1640: current_page <= 12'd1841;
            12'd1641: current_page <= 12'd310;
            12'd1642: current_page <= 12'd832;
            12'd1643: current_page <= 12'd1354;
            12'd1644: current_page <= 12'd1876;
            12'd1645: current_page <= 12'd345;
            12'd1646: current_page <= 12'd867;
            12'd1647: current_page <= 12'd1389;
            12'd1648: current_page <= 12'd1911;
            12'd1649: current_page <= 12'd380;
            12'd1650: current_page <= 12'd902;
            12'd1651: current_page <= 12'd1424;
            12'd1652: current_page <= 12'd1946;
            12'd1653: current_page <= 12'd415;
            12'd1654: current_page <= 12'd937;
            12'd1655: current_page <= 12'd1459;
            12'd1656: current_page <= 12'd1981;
            12'd1657: current_page <= 12'd450;
            12'd1658: current_page <= 12'd972;
            12'd1659: current_page <= 12'd1494;
            12'd1660: current_page <= 12'd2016;
            12'd1661: current_page <= 12'd485;
            12'd1662: current_page <= 12'd1007;
            12'd1663: current_page <= 12'd1529;
            12'd1664: current_page <= 12'd2051;
            12'd1665: current_page <= 12'd520;
            12'd1666: current_page <= 12'd1042;
            12'd1667: current_page <= 12'd1564;
            12'd1668: current_page <= 12'd33;
            12'd1669: current_page <= 12'd555;
            12'd1670: current_page <= 12'd1077;
            12'd1671: current_page <= 12'd1599;
            12'd1672: current_page <= 12'd68;
            12'd1673: current_page <= 12'd590;
            12'd1674: current_page <= 12'd1112;
            12'd1675: current_page <= 12'd1634;
            12'd1676: current_page <= 12'd103;
            12'd1677: current_page <= 12'd625;
            12'd1678: current_page <= 12'd1147;
            12'd1679: current_page <= 12'd1669;
            12'd1680: current_page <= 12'd138;
            12'd1681: current_page <= 12'd660;
            12'd1682: current_page <= 12'd1182;
            12'd1683: current_page <= 12'd1704;
            12'd1684: current_page <= 12'd173;
            12'd1685: current_page <= 12'd695;
            12'd1686: current_page <= 12'd1217;
            12'd1687: current_page <= 12'd1739;
            12'd1688: current_page <= 12'd208;
            12'd1689: current_page <= 12'd730;
            12'd1690: current_page <= 12'd1252;
            12'd1691: current_page <= 12'd1774;
            12'd1692: current_page <= 12'd243;
            12'd1693: current_page <= 12'd765;
            12'd1694: current_page <= 12'd1287;
            12'd1695: current_page <= 12'd1809;
            12'd1696: current_page <= 12'd278;
            12'd1697: current_page <= 12'd800;
            12'd1698: current_page <= 12'd1322;
            12'd1699: current_page <= 12'd1844;
            12'd1700: current_page <= 12'd313;
            12'd1701: current_page <= 12'd835;
            12'd1702: current_page <= 12'd1357;
            12'd1703: current_page <= 12'd1879;
            12'd1704: current_page <= 12'd348;
            12'd1705: current_page <= 12'd870;
            12'd1706: current_page <= 12'd1392;
            12'd1707: current_page <= 12'd1914;
            12'd1708: current_page <= 12'd383;
            12'd1709: current_page <= 12'd905;
            12'd1710: current_page <= 12'd1427;
            12'd1711: current_page <= 12'd1949;
            12'd1712: current_page <= 12'd418;
            12'd1713: current_page <= 12'd940;
            12'd1714: current_page <= 12'd1462;
            12'd1715: current_page <= 12'd1984;
            12'd1716: current_page <= 12'd453;
            12'd1717: current_page <= 12'd975;
            12'd1718: current_page <= 12'd1497;
            12'd1719: current_page <= 12'd2019;
            12'd1720: current_page <= 12'd488;
            12'd1721: current_page <= 12'd1010;
            12'd1722: current_page <= 12'd1532;
            12'd1723: current_page <= 12'd1;
            12'd1724: current_page <= 12'd523;
            12'd1725: current_page <= 12'd1045;
            12'd1726: current_page <= 12'd1567;
            12'd1727: current_page <= 12'd36;
            12'd1728: current_page <= 12'd558;
            12'd1729: current_page <= 12'd1080;
            12'd1730: current_page <= 12'd1602;
            12'd1731: current_page <= 12'd71;
            12'd1732: current_page <= 12'd593;
            12'd1733: current_page <= 12'd1115;
            12'd1734: current_page <= 12'd1637;
            12'd1735: current_page <= 12'd106;
            12'd1736: current_page <= 12'd628;
            12'd1737: current_page <= 12'd1150;
            12'd1738: current_page <= 12'd1672;
            12'd1739: current_page <= 12'd141;
            12'd1740: current_page <= 12'd663;
            12'd1741: current_page <= 12'd1185;
            12'd1742: current_page <= 12'd1707;
            12'd1743: current_page <= 12'd176;
            12'd1744: current_page <= 12'd698;
            12'd1745: current_page <= 12'd1220;
            12'd1746: current_page <= 12'd1742;
            12'd1747: current_page <= 12'd211;
            12'd1748: current_page <= 12'd733;
            12'd1749: current_page <= 12'd1255;
            12'd1750: current_page <= 12'd1777;
            12'd1751: current_page <= 12'd246;
            12'd1752: current_page <= 12'd768;
            12'd1753: current_page <= 12'd1290;
            12'd1754: current_page <= 12'd1812;
            12'd1755: current_page <= 12'd281;
            12'd1756: current_page <= 12'd803;
            12'd1757: current_page <= 12'd1325;
            12'd1758: current_page <= 12'd1847;
            12'd1759: current_page <= 12'd316;
            12'd1760: current_page <= 12'd838;
            12'd1761: current_page <= 12'd1360;
            12'd1762: current_page <= 12'd1882;
            12'd1763: current_page <= 12'd351;
            12'd1764: current_page <= 12'd873;
            12'd1765: current_page <= 12'd1395;
            12'd1766: current_page <= 12'd1917;
            12'd1767: current_page <= 12'd386;
            12'd1768: current_page <= 12'd908;
            12'd1769: current_page <= 12'd1430;
            12'd1770: current_page <= 12'd1952;
            12'd1771: current_page <= 12'd421;
            12'd1772: current_page <= 12'd943;
            12'd1773: current_page <= 12'd1465;
            12'd1774: current_page <= 12'd1987;
            12'd1775: current_page <= 12'd456;
            12'd1776: current_page <= 12'd978;
            12'd1777: current_page <= 12'd1500;
            12'd1778: current_page <= 12'd2022;
            12'd1779: current_page <= 12'd491;
            12'd1780: current_page <= 12'd1013;
            12'd1781: current_page <= 12'd1535;
            12'd1782: current_page <= 12'd4;
            12'd1783: current_page <= 12'd526;
            12'd1784: current_page <= 12'd1048;
            12'd1785: current_page <= 12'd1570;
            12'd1786: current_page <= 12'd39;
            12'd1787: current_page <= 12'd561;
            12'd1788: current_page <= 12'd1083;
            12'd1789: current_page <= 12'd1605;
            12'd1790: current_page <= 12'd74;
            12'd1791: current_page <= 12'd596;
            12'd1792: current_page <= 12'd1118;
            12'd1793: current_page <= 12'd1640;
            12'd1794: current_page <= 12'd109;
            12'd1795: current_page <= 12'd631;
            12'd1796: current_page <= 12'd1153;
            12'd1797: current_page <= 12'd1675;
            12'd1798: current_page <= 12'd144;
            12'd1799: current_page <= 12'd666;
            12'd1800: current_page <= 12'd1188;
            12'd1801: current_page <= 12'd1710;
            12'd1802: current_page <= 12'd179;
            12'd1803: current_page <= 12'd701;
            12'd1804: current_page <= 12'd1223;
            12'd1805: current_page <= 12'd1745;
            12'd1806: current_page <= 12'd214;
            12'd1807: current_page <= 12'd736;
            12'd1808: current_page <= 12'd1258;
            12'd1809: current_page <= 12'd1780;
            12'd1810: current_page <= 12'd249;
            12'd1811: current_page <= 12'd771;
            12'd1812: current_page <= 12'd1293;
            12'd1813: current_page <= 12'd1815;
            12'd1814: current_page <= 12'd284;
            12'd1815: current_page <= 12'd806;
            12'd1816: current_page <= 12'd1328;
            12'd1817: current_page <= 12'd1850;
            12'd1818: current_page <= 12'd319;
            12'd1819: current_page <= 12'd841;
            12'd1820: current_page <= 12'd1363;
            12'd1821: current_page <= 12'd1885;
            12'd1822: current_page <= 12'd354;
            12'd1823: current_page <= 12'd876;
            12'd1824: current_page <= 12'd1398;
            12'd1825: current_page <= 12'd1920;
            12'd1826: current_page <= 12'd389;
            12'd1827: current_page <= 12'd911;
            12'd1828: current_page <= 12'd1433;
            12'd1829: current_page <= 12'd1955;
            12'd1830: current_page <= 12'd424;
            12'd1831: current_page <= 12'd946;
            12'd1832: current_page <= 12'd1468;
            12'd1833: current_page <= 12'd1990;
            12'd1834: current_page <= 12'd459;
            12'd1835: current_page <= 12'd981;
            12'd1836: current_page <= 12'd1503;
            12'd1837: current_page <= 12'd2025;
            12'd1838: current_page <= 12'd494;
            12'd1839: current_page <= 12'd1016;
            12'd1840: current_page <= 12'd1538;
            12'd1841: current_page <= 12'd7;
            12'd1842: current_page <= 12'd529;
            12'd1843: current_page <= 12'd1051;
            12'd1844: current_page <= 12'd1573;
            12'd1845: current_page <= 12'd42;
            12'd1846: current_page <= 12'd564;
            12'd1847: current_page <= 12'd1086;
            12'd1848: current_page <= 12'd1608;
            12'd1849: current_page <= 12'd77;
            12'd1850: current_page <= 12'd599;
            12'd1851: current_page <= 12'd1121;
            12'd1852: current_page <= 12'd1643;
            12'd1853: current_page <= 12'd112;
            12'd1854: current_page <= 12'd634;
            12'd1855: current_page <= 12'd1156;
            12'd1856: current_page <= 12'd1678;
            12'd1857: current_page <= 12'd147;
            12'd1858: current_page <= 12'd669;
            12'd1859: current_page <= 12'd1191;
            12'd1860: current_page <= 12'd1713;
            12'd1861: current_page <= 12'd182;
            12'd1862: current_page <= 12'd704;
            12'd1863: current_page <= 12'd1226;
            12'd1864: current_page <= 12'd1748;
            12'd1865: current_page <= 12'd217;
            12'd1866: current_page <= 12'd739;
            12'd1867: current_page <= 12'd1261;
            12'd1868: current_page <= 12'd1783;
            12'd1869: current_page <= 12'd252;
            12'd1870: current_page <= 12'd774;
            12'd1871: current_page <= 12'd1296;
            12'd1872: current_page <= 12'd1818;
            12'd1873: current_page <= 12'd287;
            12'd1874: current_page <= 12'd809;
            12'd1875: current_page <= 12'd1331;
            12'd1876: current_page <= 12'd1853;
            12'd1877: current_page <= 12'd322;
            12'd1878: current_page <= 12'd844;
            12'd1879: current_page <= 12'd1366;
            12'd1880: current_page <= 12'd1888;
            12'd1881: current_page <= 12'd357;
            12'd1882: current_page <= 12'd879;
            12'd1883: current_page <= 12'd1401;
            12'd1884: current_page <= 12'd1923;
            12'd1885: current_page <= 12'd392;
            12'd1886: current_page <= 12'd914;
            12'd1887: current_page <= 12'd1436;
            12'd1888: current_page <= 12'd1958;
            12'd1889: current_page <= 12'd427;
            12'd1890: current_page <= 12'd949;
            12'd1891: current_page <= 12'd1471;
            12'd1892: current_page <= 12'd1993;
            12'd1893: current_page <= 12'd462;
            12'd1894: current_page <= 12'd984;
            12'd1895: current_page <= 12'd1506;
            12'd1896: current_page <= 12'd2028;
            12'd1897: current_page <= 12'd497;
            12'd1898: current_page <= 12'd1019;
            12'd1899: current_page <= 12'd1541;
            12'd1900: current_page <= 12'd10;
            12'd1901: current_page <= 12'd532;
            12'd1902: current_page <= 12'd1054;
            12'd1903: current_page <= 12'd1576;
            12'd1904: current_page <= 12'd45;
            12'd1905: current_page <= 12'd567;
            12'd1906: current_page <= 12'd1089;
            12'd1907: current_page <= 12'd1611;
            12'd1908: current_page <= 12'd80;
            12'd1909: current_page <= 12'd602;
            12'd1910: current_page <= 12'd1124;
            12'd1911: current_page <= 12'd1646;
            12'd1912: current_page <= 12'd115;
            12'd1913: current_page <= 12'd637;
            12'd1914: current_page <= 12'd1159;
            12'd1915: current_page <= 12'd1681;
            12'd1916: current_page <= 12'd150;
            12'd1917: current_page <= 12'd672;
            12'd1918: current_page <= 12'd1194;
            12'd1919: current_page <= 12'd1716;
            12'd1920: current_page <= 12'd185;
            12'd1921: current_page <= 12'd707;
            12'd1922: current_page <= 12'd1229;
            12'd1923: current_page <= 12'd1751;
            12'd1924: current_page <= 12'd220;
            12'd1925: current_page <= 12'd742;
            12'd1926: current_page <= 12'd1264;
            12'd1927: current_page <= 12'd1786;
            12'd1928: current_page <= 12'd255;
            12'd1929: current_page <= 12'd777;
            12'd1930: current_page <= 12'd1299;
            12'd1931: current_page <= 12'd1821;
            12'd1932: current_page <= 12'd290;
            12'd1933: current_page <= 12'd812;
            12'd1934: current_page <= 12'd1334;
            12'd1935: current_page <= 12'd1856;
            12'd1936: current_page <= 12'd325;
            12'd1937: current_page <= 12'd847;
            12'd1938: current_page <= 12'd1369;
            12'd1939: current_page <= 12'd1891;
            12'd1940: current_page <= 12'd360;
            12'd1941: current_page <= 12'd882;
            12'd1942: current_page <= 12'd1404;
            12'd1943: current_page <= 12'd1926;
            12'd1944: current_page <= 12'd395;
            12'd1945: current_page <= 12'd917;
            12'd1946: current_page <= 12'd1439;
            12'd1947: current_page <= 12'd1961;
            12'd1948: current_page <= 12'd430;
            12'd1949: current_page <= 12'd952;
            12'd1950: current_page <= 12'd1474;
            12'd1951: current_page <= 12'd1996;
            12'd1952: current_page <= 12'd465;
            12'd1953: current_page <= 12'd987;
            12'd1954: current_page <= 12'd1509;
            12'd1955: current_page <= 12'd2031;
            12'd1956: current_page <= 12'd500;
            12'd1957: current_page <= 12'd1022;
            12'd1958: current_page <= 12'd1544;
            12'd1959: current_page <= 12'd13;
            12'd1960: current_page <= 12'd535;
            12'd1961: current_page <= 12'd1057;
            12'd1962: current_page <= 12'd1579;
            12'd1963: current_page <= 12'd48;
            12'd1964: current_page <= 12'd570;
            12'd1965: current_page <= 12'd1092;
            12'd1966: current_page <= 12'd1614;
            12'd1967: current_page <= 12'd83;
            12'd1968: current_page <= 12'd605;
            12'd1969: current_page <= 12'd1127;
            12'd1970: current_page <= 12'd1649;
            12'd1971: current_page <= 12'd118;
            12'd1972: current_page <= 12'd640;
            12'd1973: current_page <= 12'd1162;
            12'd1974: current_page <= 12'd1684;
            12'd1975: current_page <= 12'd153;
            12'd1976: current_page <= 12'd675;
            12'd1977: current_page <= 12'd1197;
            12'd1978: current_page <= 12'd1719;
            12'd1979: current_page <= 12'd188;
            12'd1980: current_page <= 12'd710;
            12'd1981: current_page <= 12'd1232;
            12'd1982: current_page <= 12'd1754;
            12'd1983: current_page <= 12'd223;
            12'd1984: current_page <= 12'd745;
            12'd1985: current_page <= 12'd1267;
            12'd1986: current_page <= 12'd1789;
            12'd1987: current_page <= 12'd258;
            12'd1988: current_page <= 12'd780;
            12'd1989: current_page <= 12'd1302;
            12'd1990: current_page <= 12'd1824;
            12'd1991: current_page <= 12'd293;
            12'd1992: current_page <= 12'd815;
            12'd1993: current_page <= 12'd1337;
            12'd1994: current_page <= 12'd1859;
            12'd1995: current_page <= 12'd328;
            12'd1996: current_page <= 12'd850;
            12'd1997: current_page <= 12'd1372;
            12'd1998: current_page <= 12'd1894;
            12'd1999: current_page <= 12'd363;
            12'd2000: current_page <= 12'd885;
            12'd2001: current_page <= 12'd1407;
            12'd2002: current_page <= 12'd1929;
            12'd2003: current_page <= 12'd398;
            12'd2004: current_page <= 12'd920;
            12'd2005: current_page <= 12'd1442;
            12'd2006: current_page <= 12'd1964;
            12'd2007: current_page <= 12'd433;
            12'd2008: current_page <= 12'd955;
            12'd2009: current_page <= 12'd1477;
            12'd2010: current_page <= 12'd1999;
            12'd2011: current_page <= 12'd468;
            12'd2012: current_page <= 12'd990;
            12'd2013: current_page <= 12'd1512;
            12'd2014: current_page <= 12'd2034;
            12'd2015: current_page <= 12'd503;
            12'd2016: current_page <= 12'd1025;
            12'd2017: current_page <= 12'd1547;
            12'd2018: current_page <= 12'd16;
            12'd2019: current_page <= 12'd538;
            12'd2020: current_page <= 12'd1060;
            12'd2021: current_page <= 12'd1582;
            12'd2022: current_page <= 12'd51;
            12'd2023: current_page <= 12'd573;
            12'd2024: current_page <= 12'd1095;
            12'd2025: current_page <= 12'd1617;
            12'd2026: current_page <= 12'd86;
            12'd2027: current_page <= 12'd608;
            12'd2028: current_page <= 12'd1130;
            12'd2029: current_page <= 12'd1652;
            12'd2030: current_page <= 12'd121;
            12'd2031: current_page <= 12'd643;
            12'd2032: current_page <= 12'd1165;
            12'd2033: current_page <= 12'd1687;
            12'd2034: current_page <= 12'd156;
            12'd2035: current_page <= 12'd678;
            12'd2036: current_page <= 12'd1200;
            12'd2037: current_page <= 12'd1722;
            12'd2038: current_page <= 12'd191;
            12'd2039: current_page <= 12'd713;
            12'd2040: current_page <= 12'd1235;
            12'd2041: current_page <= 12'd1757;
            12'd2042: current_page <= 12'd226;
            12'd2043: current_page <= 12'd748;
            12'd2044: current_page <= 12'd1270;
            12'd2045: current_page <= 12'd1792;
            12'd2046: current_page <= 12'd261;
            12'd2047: current_page <= 12'd783;
            12'd2048: current_page <= 12'd1305;
            12'd2049: current_page <= 12'd1827;
            12'd2050: current_page <= 12'd296;
            12'd2051: current_page <= 12'd818;
            12'd2052: current_page <= 12'd1340;
            12'd2053: current_page <= 12'd4095;
            12'd2054: current_page <= 12'd4095;
            12'd2055: current_page <= 12'd4095;
            12'd2056: current_page <= 12'd4095;
            12'd2057: current_page <= 12'd4095;
            12'd2058: current_page <= 12'd4095;
            12'd2059: current_page <= 12'd4095;
            12'd2060: current_page <= 12'd4095;
            12'd2061: current_page <= 12'd4095;
            12'd2062: current_page <= 12'd4095;
            12'd2063: current_page <= 12'd4095;
            12'd2064: current_page <= 12'd4095;
            12'd2065: current_page <= 12'd4095;
            12'd2066: current_page <= 12'd4095;
            12'd2067: current_page <= 12'd4095;
            12'd2068: current_page <= 12'd4095;
            12'd2069: current_page <= 12'd4095;
            12'd2070: current_page <= 12'd4095;
            12'd2071: current_page <= 12'd4095;
            12'd2072: current_page <= 12'd4095;
            12'd2073: current_page <= 12'd4095;
            12'd2074: current_page <= 12'd4095;
            12'd2075: current_page <= 12'd4095;
            12'd2076: current_page <= 12'd4095;
            12'd2077: current_page <= 12'd4095;
            12'd2078: current_page <= 12'd4095;
            12'd2079: current_page <= 12'd4095;
            12'd2080: current_page <= 12'd4095;
            12'd2081: current_page <= 12'd4095;
            12'd2082: current_page <= 12'd4095;
            12'd2083: current_page <= 12'd4095;
            12'd2084: current_page <= 12'd4095;
            12'd2085: current_page <= 12'd4095;
            12'd2086: current_page <= 12'd4095;
            12'd2087: current_page <= 12'd4095;
            12'd2088: current_page <= 12'd4095;
            12'd2089: current_page <= 12'd4095;
            12'd2090: current_page <= 12'd4095;
            12'd2091: current_page <= 12'd4095;
            12'd2092: current_page <= 12'd4095;
            12'd2093: current_page <= 12'd4095;
            12'd2094: current_page <= 12'd4095;
            12'd2095: current_page <= 12'd4095;
            12'd2096: current_page <= 12'd4095;
            12'd2097: current_page <= 12'd4095;
            12'd2098: current_page <= 12'd4095;
            12'd2099: current_page <= 12'd4095;
            12'd2100: current_page <= 12'd4095;
            12'd2101: current_page <= 12'd4095;
            12'd2102: current_page <= 12'd4095;
            12'd2103: current_page <= 12'd4095;
            12'd2104: current_page <= 12'd4095;
            12'd2105: current_page <= 12'd4095;
            12'd2106: current_page <= 12'd4095;
            12'd2107: current_page <= 12'd4095;
            12'd2108: current_page <= 12'd4095;
            12'd2109: current_page <= 12'd4095;
            12'd2110: current_page <= 12'd4095;
            12'd2111: current_page <= 12'd4095;
            12'd2112: current_page <= 12'd4095;
            12'd2113: current_page <= 12'd4095;
            12'd2114: current_page <= 12'd4095;
            12'd2115: current_page <= 12'd4095;
            12'd2116: current_page <= 12'd4095;
            12'd2117: current_page <= 12'd4095;
            12'd2118: current_page <= 12'd4095;
            12'd2119: current_page <= 12'd4095;
            12'd2120: current_page <= 12'd4095;
            12'd2121: current_page <= 12'd4095;
            12'd2122: current_page <= 12'd4095;
            12'd2123: current_page <= 12'd4095;
            12'd2124: current_page <= 12'd4095;
            12'd2125: current_page <= 12'd4095;
            12'd2126: current_page <= 12'd4095;
            12'd2127: current_page <= 12'd4095;
            12'd2128: current_page <= 12'd4095;
            12'd2129: current_page <= 12'd4095;
            12'd2130: current_page <= 12'd4095;
            12'd2131: current_page <= 12'd4095;
            12'd2132: current_page <= 12'd4095;
            12'd2133: current_page <= 12'd4095;
            12'd2134: current_page <= 12'd4095;
            12'd2135: current_page <= 12'd4095;
            12'd2136: current_page <= 12'd4095;
            12'd2137: current_page <= 12'd4095;
            12'd2138: current_page <= 12'd4095;
            12'd2139: current_page <= 12'd4095;
            12'd2140: current_page <= 12'd4095;
            12'd2141: current_page <= 12'd4095;
            12'd2142: current_page <= 12'd4095;
            12'd2143: current_page <= 12'd4095;
            12'd2144: current_page <= 12'd4095;
            12'd2145: current_page <= 12'd4095;
            12'd2146: current_page <= 12'd4095;
            12'd2147: current_page <= 12'd4095;
            12'd2148: current_page <= 12'd4095;
            12'd2149: current_page <= 12'd4095;
            12'd2150: current_page <= 12'd4095;
            12'd2151: current_page <= 12'd4095;
            12'd2152: current_page <= 12'd4095;
            12'd2153: current_page <= 12'd4095;
            12'd2154: current_page <= 12'd4095;
            12'd2155: current_page <= 12'd4095;
            12'd2156: current_page <= 12'd4095;
            12'd2157: current_page <= 12'd4095;
            12'd2158: current_page <= 12'd4095;
            12'd2159: current_page <= 12'd4095;
            12'd2160: current_page <= 12'd4095;
            12'd2161: current_page <= 12'd4095;
            12'd2162: current_page <= 12'd4095;
            12'd2163: current_page <= 12'd4095;
            12'd2164: current_page <= 12'd4095;
            12'd2165: current_page <= 12'd4095;
            12'd2166: current_page <= 12'd4095;
            12'd2167: current_page <= 12'd4095;
            12'd2168: current_page <= 12'd4095;
            12'd2169: current_page <= 12'd4095;
            12'd2170: current_page <= 12'd4095;
            12'd2171: current_page <= 12'd4095;
            12'd2172: current_page <= 12'd4095;
            12'd2173: current_page <= 12'd4095;
            12'd2174: current_page <= 12'd4095;
            12'd2175: current_page <= 12'd4095;
            12'd2176: current_page <= 12'd4095;
            12'd2177: current_page <= 12'd4095;
            12'd2178: current_page <= 12'd4095;
            12'd2179: current_page <= 12'd4095;
            12'd2180: current_page <= 12'd4095;
            12'd2181: current_page <= 12'd4095;
            12'd2182: current_page <= 12'd4095;
            12'd2183: current_page <= 12'd4095;
            12'd2184: current_page <= 12'd4095;
            12'd2185: current_page <= 12'd4095;
            12'd2186: current_page <= 12'd4095;
            12'd2187: current_page <= 12'd4095;
            12'd2188: current_page <= 12'd4095;
            12'd2189: current_page <= 12'd4095;
            12'd2190: current_page <= 12'd4095;
            12'd2191: current_page <= 12'd4095;
            12'd2192: current_page <= 12'd4095;
            12'd2193: current_page <= 12'd4095;
            12'd2194: current_page <= 12'd4095;
            12'd2195: current_page <= 12'd4095;
            12'd2196: current_page <= 12'd4095;
            12'd2197: current_page <= 12'd4095;
            12'd2198: current_page <= 12'd4095;
            12'd2199: current_page <= 12'd4095;
            12'd2200: current_page <= 12'd4095;
            12'd2201: current_page <= 12'd4095;
            12'd2202: current_page <= 12'd4095;
            12'd2203: current_page <= 12'd4095;
            12'd2204: current_page <= 12'd4095;
            12'd2205: current_page <= 12'd4095;
            12'd2206: current_page <= 12'd4095;
            12'd2207: current_page <= 12'd4095;
            12'd2208: current_page <= 12'd4095;
            12'd2209: current_page <= 12'd4095;
            12'd2210: current_page <= 12'd4095;
            12'd2211: current_page <= 12'd4095;
            12'd2212: current_page <= 12'd4095;
            12'd2213: current_page <= 12'd4095;
            12'd2214: current_page <= 12'd4095;
            12'd2215: current_page <= 12'd4095;
            12'd2216: current_page <= 12'd4095;
            12'd2217: current_page <= 12'd4095;
            12'd2218: current_page <= 12'd4095;
            12'd2219: current_page <= 12'd4095;
            12'd2220: current_page <= 12'd4095;
            12'd2221: current_page <= 12'd4095;
            12'd2222: current_page <= 12'd4095;
            12'd2223: current_page <= 12'd4095;
            12'd2224: current_page <= 12'd4095;
            12'd2225: current_page <= 12'd4095;
            12'd2226: current_page <= 12'd4095;
            12'd2227: current_page <= 12'd4095;
            12'd2228: current_page <= 12'd4095;
            12'd2229: current_page <= 12'd4095;
            12'd2230: current_page <= 12'd4095;
            12'd2231: current_page <= 12'd4095;
            12'd2232: current_page <= 12'd4095;
            12'd2233: current_page <= 12'd4095;
            12'd2234: current_page <= 12'd4095;
            12'd2235: current_page <= 12'd4095;
            12'd2236: current_page <= 12'd4095;
            12'd2237: current_page <= 12'd4095;
            12'd2238: current_page <= 12'd4095;
            12'd2239: current_page <= 12'd4095;
            12'd2240: current_page <= 12'd4095;
            12'd2241: current_page <= 12'd4095;
            12'd2242: current_page <= 12'd4095;
            12'd2243: current_page <= 12'd4095;
            12'd2244: current_page <= 12'd4095;
            12'd2245: current_page <= 12'd4095;
            12'd2246: current_page <= 12'd4095;
            12'd2247: current_page <= 12'd4095;
            12'd2248: current_page <= 12'd4095;
            12'd2249: current_page <= 12'd4095;
            12'd2250: current_page <= 12'd4095;
            12'd2251: current_page <= 12'd4095;
            12'd2252: current_page <= 12'd4095;
            12'd2253: current_page <= 12'd4095;
            12'd2254: current_page <= 12'd4095;
            12'd2255: current_page <= 12'd4095;
            12'd2256: current_page <= 12'd4095;
            12'd2257: current_page <= 12'd4095;
            12'd2258: current_page <= 12'd4095;
            12'd2259: current_page <= 12'd4095;
            12'd2260: current_page <= 12'd4095;
            12'd2261: current_page <= 12'd4095;
            12'd2262: current_page <= 12'd4095;
            12'd2263: current_page <= 12'd4095;
            12'd2264: current_page <= 12'd4095;
            12'd2265: current_page <= 12'd4095;
            12'd2266: current_page <= 12'd4095;
            12'd2267: current_page <= 12'd4095;
            12'd2268: current_page <= 12'd4095;
            12'd2269: current_page <= 12'd4095;
            12'd2270: current_page <= 12'd4095;
            12'd2271: current_page <= 12'd4095;
            12'd2272: current_page <= 12'd4095;
            12'd2273: current_page <= 12'd4095;
            12'd2274: current_page <= 12'd4095;
            12'd2275: current_page <= 12'd4095;
            12'd2276: current_page <= 12'd4095;
            12'd2277: current_page <= 12'd4095;
            12'd2278: current_page <= 12'd4095;
            12'd2279: current_page <= 12'd4095;
            12'd2280: current_page <= 12'd4095;
            12'd2281: current_page <= 12'd4095;
            12'd2282: current_page <= 12'd4095;
            12'd2283: current_page <= 12'd4095;
            12'd2284: current_page <= 12'd4095;
            12'd2285: current_page <= 12'd4095;
            12'd2286: current_page <= 12'd4095;
            12'd2287: current_page <= 12'd4095;
            12'd2288: current_page <= 12'd4095;
            12'd2289: current_page <= 12'd4095;
            12'd2290: current_page <= 12'd4095;
            12'd2291: current_page <= 12'd4095;
            12'd2292: current_page <= 12'd4095;
            12'd2293: current_page <= 12'd4095;
            12'd2294: current_page <= 12'd4095;
            12'd2295: current_page <= 12'd4095;
            12'd2296: current_page <= 12'd4095;
            12'd2297: current_page <= 12'd4095;
            12'd2298: current_page <= 12'd4095;
            12'd2299: current_page <= 12'd4095;
            12'd2300: current_page <= 12'd4095;
            12'd2301: current_page <= 12'd4095;
            12'd2302: current_page <= 12'd4095;
            12'd2303: current_page <= 12'd4095;
            12'd2304: current_page <= 12'd4095;
            12'd2305: current_page <= 12'd4095;
            12'd2306: current_page <= 12'd4095;
            12'd2307: current_page <= 12'd4095;
            12'd2308: current_page <= 12'd4095;
            12'd2309: current_page <= 12'd4095;
            12'd2310: current_page <= 12'd4095;
            12'd2311: current_page <= 12'd4095;
            12'd2312: current_page <= 12'd4095;
            12'd2313: current_page <= 12'd4095;
            12'd2314: current_page <= 12'd4095;
            12'd2315: current_page <= 12'd4095;
            12'd2316: current_page <= 12'd4095;
            12'd2317: current_page <= 12'd4095;
            12'd2318: current_page <= 12'd4095;
            12'd2319: current_page <= 12'd4095;
            12'd2320: current_page <= 12'd4095;
            12'd2321: current_page <= 12'd4095;
            12'd2322: current_page <= 12'd4095;
            12'd2323: current_page <= 12'd4095;
            12'd2324: current_page <= 12'd4095;
            12'd2325: current_page <= 12'd4095;
            12'd2326: current_page <= 12'd4095;
            12'd2327: current_page <= 12'd4095;
            12'd2328: current_page <= 12'd4095;
            12'd2329: current_page <= 12'd4095;
            12'd2330: current_page <= 12'd4095;
            12'd2331: current_page <= 12'd4095;
            12'd2332: current_page <= 12'd4095;
            12'd2333: current_page <= 12'd4095;
            12'd2334: current_page <= 12'd4095;
            12'd2335: current_page <= 12'd4095;
            12'd2336: current_page <= 12'd4095;
            12'd2337: current_page <= 12'd4095;
            12'd2338: current_page <= 12'd4095;
            12'd2339: current_page <= 12'd4095;
            12'd2340: current_page <= 12'd4095;
            12'd2341: current_page <= 12'd4095;
            12'd2342: current_page <= 12'd4095;
            12'd2343: current_page <= 12'd4095;
            12'd2344: current_page <= 12'd4095;
            12'd2345: current_page <= 12'd4095;
            12'd2346: current_page <= 12'd4095;
            12'd2347: current_page <= 12'd4095;
            12'd2348: current_page <= 12'd4095;
            12'd2349: current_page <= 12'd4095;
            12'd2350: current_page <= 12'd4095;
            12'd2351: current_page <= 12'd4095;
            12'd2352: current_page <= 12'd4095;
            12'd2353: current_page <= 12'd4095;
            12'd2354: current_page <= 12'd4095;
            12'd2355: current_page <= 12'd4095;
            12'd2356: current_page <= 12'd4095;
            12'd2357: current_page <= 12'd4095;
            12'd2358: current_page <= 12'd4095;
            12'd2359: current_page <= 12'd4095;
            12'd2360: current_page <= 12'd4095;
            12'd2361: current_page <= 12'd4095;
            12'd2362: current_page <= 12'd4095;
            12'd2363: current_page <= 12'd4095;
            12'd2364: current_page <= 12'd4095;
            12'd2365: current_page <= 12'd4095;
            12'd2366: current_page <= 12'd4095;
            12'd2367: current_page <= 12'd4095;
            12'd2368: current_page <= 12'd4095;
            12'd2369: current_page <= 12'd4095;
            12'd2370: current_page <= 12'd4095;
            12'd2371: current_page <= 12'd4095;
            12'd2372: current_page <= 12'd4095;
            12'd2373: current_page <= 12'd4095;
            12'd2374: current_page <= 12'd4095;
            12'd2375: current_page <= 12'd4095;
            12'd2376: current_page <= 12'd4095;
            12'd2377: current_page <= 12'd4095;
            12'd2378: current_page <= 12'd4095;
            12'd2379: current_page <= 12'd4095;
            12'd2380: current_page <= 12'd4095;
            12'd2381: current_page <= 12'd4095;
            12'd2382: current_page <= 12'd4095;
            12'd2383: current_page <= 12'd4095;
            12'd2384: current_page <= 12'd4095;
            12'd2385: current_page <= 12'd4095;
            12'd2386: current_page <= 12'd4095;
            12'd2387: current_page <= 12'd4095;
            12'd2388: current_page <= 12'd4095;
            12'd2389: current_page <= 12'd4095;
            12'd2390: current_page <= 12'd4095;
            12'd2391: current_page <= 12'd4095;
            12'd2392: current_page <= 12'd4095;
            12'd2393: current_page <= 12'd4095;
            12'd2394: current_page <= 12'd4095;
            12'd2395: current_page <= 12'd4095;
            12'd2396: current_page <= 12'd4095;
            12'd2397: current_page <= 12'd4095;
            12'd2398: current_page <= 12'd4095;
            12'd2399: current_page <= 12'd4095;
            12'd2400: current_page <= 12'd4095;
            12'd2401: current_page <= 12'd4095;
            12'd2402: current_page <= 12'd4095;
            12'd2403: current_page <= 12'd4095;
            12'd2404: current_page <= 12'd4095;
            12'd2405: current_page <= 12'd4095;
            12'd2406: current_page <= 12'd4095;
            12'd2407: current_page <= 12'd4095;
            12'd2408: current_page <= 12'd4095;
            12'd2409: current_page <= 12'd4095;
            12'd2410: current_page <= 12'd4095;
            12'd2411: current_page <= 12'd4095;
            12'd2412: current_page <= 12'd4095;
            12'd2413: current_page <= 12'd4095;
            12'd2414: current_page <= 12'd4095;
            12'd2415: current_page <= 12'd4095;
            12'd2416: current_page <= 12'd4095;
            12'd2417: current_page <= 12'd4095;
            12'd2418: current_page <= 12'd4095;
            12'd2419: current_page <= 12'd4095;
            12'd2420: current_page <= 12'd4095;
            12'd2421: current_page <= 12'd4095;
            12'd2422: current_page <= 12'd4095;
            12'd2423: current_page <= 12'd4095;
            12'd2424: current_page <= 12'd4095;
            12'd2425: current_page <= 12'd4095;
            12'd2426: current_page <= 12'd4095;
            12'd2427: current_page <= 12'd4095;
            12'd2428: current_page <= 12'd4095;
            12'd2429: current_page <= 12'd4095;
            12'd2430: current_page <= 12'd4095;
            12'd2431: current_page <= 12'd4095;
            12'd2432: current_page <= 12'd4095;
            12'd2433: current_page <= 12'd4095;
            12'd2434: current_page <= 12'd4095;
            12'd2435: current_page <= 12'd4095;
            12'd2436: current_page <= 12'd4095;
            12'd2437: current_page <= 12'd4095;
            12'd2438: current_page <= 12'd4095;
            12'd2439: current_page <= 12'd4095;
            12'd2440: current_page <= 12'd4095;
            12'd2441: current_page <= 12'd4095;
            12'd2442: current_page <= 12'd4095;
            12'd2443: current_page <= 12'd4095;
            12'd2444: current_page <= 12'd4095;
            12'd2445: current_page <= 12'd4095;
            12'd2446: current_page <= 12'd4095;
            12'd2447: current_page <= 12'd4095;
            12'd2448: current_page <= 12'd4095;
            12'd2449: current_page <= 12'd4095;
            12'd2450: current_page <= 12'd4095;
            12'd2451: current_page <= 12'd4095;
            12'd2452: current_page <= 12'd4095;
            12'd2453: current_page <= 12'd4095;
            12'd2454: current_page <= 12'd4095;
            12'd2455: current_page <= 12'd4095;
            12'd2456: current_page <= 12'd4095;
            12'd2457: current_page <= 12'd4095;
            12'd2458: current_page <= 12'd4095;
            12'd2459: current_page <= 12'd4095;
            12'd2460: current_page <= 12'd4095;
            12'd2461: current_page <= 12'd4095;
            12'd2462: current_page <= 12'd4095;
            12'd2463: current_page <= 12'd4095;
            12'd2464: current_page <= 12'd4095;
            12'd2465: current_page <= 12'd4095;
            12'd2466: current_page <= 12'd4095;
            12'd2467: current_page <= 12'd4095;
            12'd2468: current_page <= 12'd4095;
            12'd2469: current_page <= 12'd4095;
            12'd2470: current_page <= 12'd4095;
            12'd2471: current_page <= 12'd4095;
            12'd2472: current_page <= 12'd4095;
            12'd2473: current_page <= 12'd4095;
            12'd2474: current_page <= 12'd4095;
            12'd2475: current_page <= 12'd4095;
            12'd2476: current_page <= 12'd4095;
            12'd2477: current_page <= 12'd4095;
            12'd2478: current_page <= 12'd4095;
            12'd2479: current_page <= 12'd4095;
            12'd2480: current_page <= 12'd4095;
            12'd2481: current_page <= 12'd4095;
            12'd2482: current_page <= 12'd4095;
            12'd2483: current_page <= 12'd4095;
            12'd2484: current_page <= 12'd4095;
            12'd2485: current_page <= 12'd4095;
            12'd2486: current_page <= 12'd4095;
            12'd2487: current_page <= 12'd4095;
            12'd2488: current_page <= 12'd4095;
            12'd2489: current_page <= 12'd4095;
            12'd2490: current_page <= 12'd4095;
            12'd2491: current_page <= 12'd4095;
            12'd2492: current_page <= 12'd4095;
            12'd2493: current_page <= 12'd4095;
            12'd2494: current_page <= 12'd4095;
            12'd2495: current_page <= 12'd4095;
            12'd2496: current_page <= 12'd4095;
            12'd2497: current_page <= 12'd4095;
            12'd2498: current_page <= 12'd4095;
            12'd2499: current_page <= 12'd4095;
            12'd2500: current_page <= 12'd4095;
            12'd2501: current_page <= 12'd4095;
            12'd2502: current_page <= 12'd4095;
            12'd2503: current_page <= 12'd4095;
            12'd2504: current_page <= 12'd4095;
            12'd2505: current_page <= 12'd4095;
            12'd2506: current_page <= 12'd4095;
            12'd2507: current_page <= 12'd4095;
            12'd2508: current_page <= 12'd4095;
            12'd2509: current_page <= 12'd4095;
            12'd2510: current_page <= 12'd4095;
            12'd2511: current_page <= 12'd4095;
            12'd2512: current_page <= 12'd4095;
            12'd2513: current_page <= 12'd4095;
            12'd2514: current_page <= 12'd4095;
            12'd2515: current_page <= 12'd4095;
            12'd2516: current_page <= 12'd4095;
            12'd2517: current_page <= 12'd4095;
            12'd2518: current_page <= 12'd4095;
            12'd2519: current_page <= 12'd4095;
            12'd2520: current_page <= 12'd4095;
            12'd2521: current_page <= 12'd4095;
            12'd2522: current_page <= 12'd4095;
            12'd2523: current_page <= 12'd4095;
            12'd2524: current_page <= 12'd4095;
            12'd2525: current_page <= 12'd4095;
            12'd2526: current_page <= 12'd4095;
            12'd2527: current_page <= 12'd4095;
            12'd2528: current_page <= 12'd4095;
            12'd2529: current_page <= 12'd4095;
            12'd2530: current_page <= 12'd4095;
            12'd2531: current_page <= 12'd4095;
            12'd2532: current_page <= 12'd4095;
            12'd2533: current_page <= 12'd4095;
            12'd2534: current_page <= 12'd4095;
            12'd2535: current_page <= 12'd4095;
            12'd2536: current_page <= 12'd4095;
            12'd2537: current_page <= 12'd4095;
            12'd2538: current_page <= 12'd4095;
            12'd2539: current_page <= 12'd4095;
            12'd2540: current_page <= 12'd4095;
            12'd2541: current_page <= 12'd4095;
            12'd2542: current_page <= 12'd4095;
            12'd2543: current_page <= 12'd4095;
            12'd2544: current_page <= 12'd4095;
            12'd2545: current_page <= 12'd4095;
            12'd2546: current_page <= 12'd4095;
            12'd2547: current_page <= 12'd4095;
            12'd2548: current_page <= 12'd4095;
            12'd2549: current_page <= 12'd4095;
            12'd2550: current_page <= 12'd4095;
            12'd2551: current_page <= 12'd4095;
            12'd2552: current_page <= 12'd4095;
            12'd2553: current_page <= 12'd4095;
            12'd2554: current_page <= 12'd4095;
            12'd2555: current_page <= 12'd4095;
            12'd2556: current_page <= 12'd4095;
            12'd2557: current_page <= 12'd4095;
            12'd2558: current_page <= 12'd4095;
            12'd2559: current_page <= 12'd4095;
            12'd2560: current_page <= 12'd4095;
            12'd2561: current_page <= 12'd4095;
            12'd2562: current_page <= 12'd4095;
            12'd2563: current_page <= 12'd4095;
            12'd2564: current_page <= 12'd4095;
            12'd2565: current_page <= 12'd4095;
            12'd2566: current_page <= 12'd4095;
            12'd2567: current_page <= 12'd4095;
            12'd2568: current_page <= 12'd4095;
            12'd2569: current_page <= 12'd4095;
            12'd2570: current_page <= 12'd4095;
            12'd2571: current_page <= 12'd4095;
            12'd2572: current_page <= 12'd4095;
            12'd2573: current_page <= 12'd4095;
            12'd2574: current_page <= 12'd4095;
            12'd2575: current_page <= 12'd4095;
            12'd2576: current_page <= 12'd4095;
            12'd2577: current_page <= 12'd4095;
            12'd2578: current_page <= 12'd4095;
            12'd2579: current_page <= 12'd4095;
            12'd2580: current_page <= 12'd4095;
            12'd2581: current_page <= 12'd4095;
            12'd2582: current_page <= 12'd4095;
            12'd2583: current_page <= 12'd4095;
            12'd2584: current_page <= 12'd4095;
            12'd2585: current_page <= 12'd4095;
            12'd2586: current_page <= 12'd4095;
            12'd2587: current_page <= 12'd4095;
            12'd2588: current_page <= 12'd4095;
            12'd2589: current_page <= 12'd4095;
            12'd2590: current_page <= 12'd4095;
            12'd2591: current_page <= 12'd4095;
            12'd2592: current_page <= 12'd4095;
            12'd2593: current_page <= 12'd4095;
            12'd2594: current_page <= 12'd4095;
            12'd2595: current_page <= 12'd4095;
            12'd2596: current_page <= 12'd4095;
            12'd2597: current_page <= 12'd4095;
            12'd2598: current_page <= 12'd4095;
            12'd2599: current_page <= 12'd4095;
            12'd2600: current_page <= 12'd4095;
            12'd2601: current_page <= 12'd4095;
            12'd2602: current_page <= 12'd4095;
            12'd2603: current_page <= 12'd4095;
            12'd2604: current_page <= 12'd4095;
            12'd2605: current_page <= 12'd4095;
            12'd2606: current_page <= 12'd4095;
            12'd2607: current_page <= 12'd4095;
            12'd2608: current_page <= 12'd4095;
            12'd2609: current_page <= 12'd4095;
            12'd2610: current_page <= 12'd4095;
            12'd2611: current_page <= 12'd4095;
            12'd2612: current_page <= 12'd4095;
            12'd2613: current_page <= 12'd4095;
            12'd2614: current_page <= 12'd4095;
            12'd2615: current_page <= 12'd4095;
            12'd2616: current_page <= 12'd4095;
            12'd2617: current_page <= 12'd4095;
            12'd2618: current_page <= 12'd4095;
            12'd2619: current_page <= 12'd4095;
            12'd2620: current_page <= 12'd4095;
            12'd2621: current_page <= 12'd4095;
            12'd2622: current_page <= 12'd4095;
            12'd2623: current_page <= 12'd4095;
            12'd2624: current_page <= 12'd4095;
            12'd2625: current_page <= 12'd4095;
            12'd2626: current_page <= 12'd4095;
            12'd2627: current_page <= 12'd4095;
            12'd2628: current_page <= 12'd4095;
            12'd2629: current_page <= 12'd4095;
            12'd2630: current_page <= 12'd4095;
            12'd2631: current_page <= 12'd4095;
            12'd2632: current_page <= 12'd4095;
            12'd2633: current_page <= 12'd4095;
            12'd2634: current_page <= 12'd4095;
            12'd2635: current_page <= 12'd4095;
            12'd2636: current_page <= 12'd4095;
            12'd2637: current_page <= 12'd4095;
            12'd2638: current_page <= 12'd4095;
            12'd2639: current_page <= 12'd4095;
            12'd2640: current_page <= 12'd4095;
            12'd2641: current_page <= 12'd4095;
            12'd2642: current_page <= 12'd4095;
            12'd2643: current_page <= 12'd4095;
            12'd2644: current_page <= 12'd4095;
            12'd2645: current_page <= 12'd4095;
            12'd2646: current_page <= 12'd4095;
            12'd2647: current_page <= 12'd4095;
            12'd2648: current_page <= 12'd4095;
            12'd2649: current_page <= 12'd4095;
            12'd2650: current_page <= 12'd4095;
            12'd2651: current_page <= 12'd4095;
            12'd2652: current_page <= 12'd4095;
            12'd2653: current_page <= 12'd4095;
            12'd2654: current_page <= 12'd4095;
            12'd2655: current_page <= 12'd4095;
            12'd2656: current_page <= 12'd4095;
            12'd2657: current_page <= 12'd4095;
            12'd2658: current_page <= 12'd4095;
            12'd2659: current_page <= 12'd4095;
            12'd2660: current_page <= 12'd4095;
            12'd2661: current_page <= 12'd4095;
            12'd2662: current_page <= 12'd4095;
            12'd2663: current_page <= 12'd4095;
            12'd2664: current_page <= 12'd4095;
            12'd2665: current_page <= 12'd4095;
            12'd2666: current_page <= 12'd4095;
            12'd2667: current_page <= 12'd4095;
            12'd2668: current_page <= 12'd4095;
            12'd2669: current_page <= 12'd4095;
            12'd2670: current_page <= 12'd4095;
            12'd2671: current_page <= 12'd4095;
            12'd2672: current_page <= 12'd4095;
            12'd2673: current_page <= 12'd4095;
            12'd2674: current_page <= 12'd4095;
            12'd2675: current_page <= 12'd4095;
            12'd2676: current_page <= 12'd4095;
            12'd2677: current_page <= 12'd4095;
            12'd2678: current_page <= 12'd4095;
            12'd2679: current_page <= 12'd4095;
            12'd2680: current_page <= 12'd4095;
            12'd2681: current_page <= 12'd4095;
            12'd2682: current_page <= 12'd4095;
            12'd2683: current_page <= 12'd4095;
            12'd2684: current_page <= 12'd4095;
            12'd2685: current_page <= 12'd4095;
            12'd2686: current_page <= 12'd4095;
            12'd2687: current_page <= 12'd4095;
            12'd2688: current_page <= 12'd4095;
            12'd2689: current_page <= 12'd4095;
            12'd2690: current_page <= 12'd4095;
            12'd2691: current_page <= 12'd4095;
            12'd2692: current_page <= 12'd4095;
            12'd2693: current_page <= 12'd4095;
            12'd2694: current_page <= 12'd4095;
            12'd2695: current_page <= 12'd4095;
            12'd2696: current_page <= 12'd4095;
            12'd2697: current_page <= 12'd4095;
            12'd2698: current_page <= 12'd4095;
            12'd2699: current_page <= 12'd4095;
            12'd2700: current_page <= 12'd4095;
            12'd2701: current_page <= 12'd4095;
            12'd2702: current_page <= 12'd4095;
            12'd2703: current_page <= 12'd4095;
            12'd2704: current_page <= 12'd4095;
            12'd2705: current_page <= 12'd4095;
            12'd2706: current_page <= 12'd4095;
            12'd2707: current_page <= 12'd4095;
            12'd2708: current_page <= 12'd4095;
            12'd2709: current_page <= 12'd4095;
            12'd2710: current_page <= 12'd4095;
            12'd2711: current_page <= 12'd4095;
            12'd2712: current_page <= 12'd4095;
            12'd2713: current_page <= 12'd4095;
            12'd2714: current_page <= 12'd4095;
            12'd2715: current_page <= 12'd4095;
            12'd2716: current_page <= 12'd4095;
            12'd2717: current_page <= 12'd4095;
            12'd2718: current_page <= 12'd4095;
            12'd2719: current_page <= 12'd4095;
            12'd2720: current_page <= 12'd4095;
            12'd2721: current_page <= 12'd4095;
            12'd2722: current_page <= 12'd4095;
            12'd2723: current_page <= 12'd4095;
            12'd2724: current_page <= 12'd4095;
            12'd2725: current_page <= 12'd4095;
            12'd2726: current_page <= 12'd4095;
            12'd2727: current_page <= 12'd4095;
            12'd2728: current_page <= 12'd4095;
            12'd2729: current_page <= 12'd4095;
            12'd2730: current_page <= 12'd4095;
            12'd2731: current_page <= 12'd4095;
            12'd2732: current_page <= 12'd4095;
            12'd2733: current_page <= 12'd4095;
            12'd2734: current_page <= 12'd4095;
            12'd2735: current_page <= 12'd4095;
            12'd2736: current_page <= 12'd4095;
            12'd2737: current_page <= 12'd4095;
            12'd2738: current_page <= 12'd4095;
            12'd2739: current_page <= 12'd4095;
            12'd2740: current_page <= 12'd4095;
            12'd2741: current_page <= 12'd4095;
            12'd2742: current_page <= 12'd4095;
            12'd2743: current_page <= 12'd4095;
            12'd2744: current_page <= 12'd4095;
            12'd2745: current_page <= 12'd4095;
            12'd2746: current_page <= 12'd4095;
            12'd2747: current_page <= 12'd4095;
            12'd2748: current_page <= 12'd4095;
            12'd2749: current_page <= 12'd4095;
            12'd2750: current_page <= 12'd4095;
            12'd2751: current_page <= 12'd4095;
            12'd2752: current_page <= 12'd4095;
            12'd2753: current_page <= 12'd4095;
            12'd2754: current_page <= 12'd4095;
            12'd2755: current_page <= 12'd4095;
            12'd2756: current_page <= 12'd4095;
            12'd2757: current_page <= 12'd4095;
            12'd2758: current_page <= 12'd4095;
            12'd2759: current_page <= 12'd4095;
            12'd2760: current_page <= 12'd4095;
            12'd2761: current_page <= 12'd4095;
            12'd2762: current_page <= 12'd4095;
            12'd2763: current_page <= 12'd4095;
            12'd2764: current_page <= 12'd4095;
            12'd2765: current_page <= 12'd4095;
            12'd2766: current_page <= 12'd4095;
            12'd2767: current_page <= 12'd4095;
            12'd2768: current_page <= 12'd4095;
            12'd2769: current_page <= 12'd4095;
            12'd2770: current_page <= 12'd4095;
            12'd2771: current_page <= 12'd4095;
            12'd2772: current_page <= 12'd4095;
            12'd2773: current_page <= 12'd4095;
            12'd2774: current_page <= 12'd4095;
            12'd2775: current_page <= 12'd4095;
            12'd2776: current_page <= 12'd4095;
            12'd2777: current_page <= 12'd4095;
            12'd2778: current_page <= 12'd4095;
            12'd2779: current_page <= 12'd4095;
            12'd2780: current_page <= 12'd4095;
            12'd2781: current_page <= 12'd4095;
            12'd2782: current_page <= 12'd4095;
            12'd2783: current_page <= 12'd4095;
            12'd2784: current_page <= 12'd4095;
            12'd2785: current_page <= 12'd4095;
            12'd2786: current_page <= 12'd4095;
            12'd2787: current_page <= 12'd4095;
            12'd2788: current_page <= 12'd4095;
            12'd2789: current_page <= 12'd4095;
            12'd2790: current_page <= 12'd4095;
            12'd2791: current_page <= 12'd4095;
            12'd2792: current_page <= 12'd4095;
            12'd2793: current_page <= 12'd4095;
            12'd2794: current_page <= 12'd4095;
            12'd2795: current_page <= 12'd4095;
            12'd2796: current_page <= 12'd4095;
            12'd2797: current_page <= 12'd4095;
            12'd2798: current_page <= 12'd4095;
            12'd2799: current_page <= 12'd4095;
            12'd2800: current_page <= 12'd4095;
            12'd2801: current_page <= 12'd4095;
            12'd2802: current_page <= 12'd4095;
            12'd2803: current_page <= 12'd4095;
            12'd2804: current_page <= 12'd4095;
            12'd2805: current_page <= 12'd4095;
            12'd2806: current_page <= 12'd4095;
            12'd2807: current_page <= 12'd4095;
            12'd2808: current_page <= 12'd4095;
            12'd2809: current_page <= 12'd4095;
            12'd2810: current_page <= 12'd4095;
            12'd2811: current_page <= 12'd4095;
            12'd2812: current_page <= 12'd4095;
            12'd2813: current_page <= 12'd4095;
            12'd2814: current_page <= 12'd4095;
            12'd2815: current_page <= 12'd4095;
            12'd2816: current_page <= 12'd4095;
            12'd2817: current_page <= 12'd4095;
            12'd2818: current_page <= 12'd4095;
            12'd2819: current_page <= 12'd4095;
            12'd2820: current_page <= 12'd4095;
            12'd2821: current_page <= 12'd4095;
            12'd2822: current_page <= 12'd4095;
            12'd2823: current_page <= 12'd4095;
            12'd2824: current_page <= 12'd4095;
            12'd2825: current_page <= 12'd4095;
            12'd2826: current_page <= 12'd4095;
            12'd2827: current_page <= 12'd4095;
            12'd2828: current_page <= 12'd4095;
            12'd2829: current_page <= 12'd4095;
            12'd2830: current_page <= 12'd4095;
            12'd2831: current_page <= 12'd4095;
            12'd2832: current_page <= 12'd4095;
            12'd2833: current_page <= 12'd4095;
            12'd2834: current_page <= 12'd4095;
            12'd2835: current_page <= 12'd4095;
            12'd2836: current_page <= 12'd4095;
            12'd2837: current_page <= 12'd4095;
            12'd2838: current_page <= 12'd4095;
            12'd2839: current_page <= 12'd4095;
            12'd2840: current_page <= 12'd4095;
            12'd2841: current_page <= 12'd4095;
            12'd2842: current_page <= 12'd4095;
            12'd2843: current_page <= 12'd4095;
            12'd2844: current_page <= 12'd4095;
            12'd2845: current_page <= 12'd4095;
            12'd2846: current_page <= 12'd4095;
            12'd2847: current_page <= 12'd4095;
            12'd2848: current_page <= 12'd4095;
            12'd2849: current_page <= 12'd4095;
            12'd2850: current_page <= 12'd4095;
            12'd2851: current_page <= 12'd4095;
            12'd2852: current_page <= 12'd4095;
            12'd2853: current_page <= 12'd4095;
            12'd2854: current_page <= 12'd4095;
            12'd2855: current_page <= 12'd4095;
            12'd2856: current_page <= 12'd4095;
            12'd2857: current_page <= 12'd4095;
            12'd2858: current_page <= 12'd4095;
            12'd2859: current_page <= 12'd4095;
            12'd2860: current_page <= 12'd4095;
            12'd2861: current_page <= 12'd4095;
            12'd2862: current_page <= 12'd4095;
            12'd2863: current_page <= 12'd4095;
            12'd2864: current_page <= 12'd4095;
            12'd2865: current_page <= 12'd4095;
            12'd2866: current_page <= 12'd4095;
            12'd2867: current_page <= 12'd4095;
            12'd2868: current_page <= 12'd4095;
            12'd2869: current_page <= 12'd4095;
            12'd2870: current_page <= 12'd4095;
            12'd2871: current_page <= 12'd4095;
            12'd2872: current_page <= 12'd4095;
            12'd2873: current_page <= 12'd4095;
            12'd2874: current_page <= 12'd4095;
            12'd2875: current_page <= 12'd4095;
            12'd2876: current_page <= 12'd4095;
            12'd2877: current_page <= 12'd4095;
            12'd2878: current_page <= 12'd4095;
            12'd2879: current_page <= 12'd4095;
            12'd2880: current_page <= 12'd4095;
            12'd2881: current_page <= 12'd4095;
            12'd2882: current_page <= 12'd4095;
            12'd2883: current_page <= 12'd4095;
            12'd2884: current_page <= 12'd4095;
            12'd2885: current_page <= 12'd4095;
            12'd2886: current_page <= 12'd4095;
            12'd2887: current_page <= 12'd4095;
            12'd2888: current_page <= 12'd4095;
            12'd2889: current_page <= 12'd4095;
            12'd2890: current_page <= 12'd4095;
            12'd2891: current_page <= 12'd4095;
            12'd2892: current_page <= 12'd4095;
            12'd2893: current_page <= 12'd4095;
            12'd2894: current_page <= 12'd4095;
            12'd2895: current_page <= 12'd4095;
            12'd2896: current_page <= 12'd4095;
            12'd2897: current_page <= 12'd4095;
            12'd2898: current_page <= 12'd4095;
            12'd2899: current_page <= 12'd4095;
            12'd2900: current_page <= 12'd4095;
            12'd2901: current_page <= 12'd4095;
            12'd2902: current_page <= 12'd4095;
            12'd2903: current_page <= 12'd4095;
            12'd2904: current_page <= 12'd4095;
            12'd2905: current_page <= 12'd4095;
            12'd2906: current_page <= 12'd4095;
            12'd2907: current_page <= 12'd4095;
            12'd2908: current_page <= 12'd4095;
            12'd2909: current_page <= 12'd4095;
            12'd2910: current_page <= 12'd4095;
            12'd2911: current_page <= 12'd4095;
            12'd2912: current_page <= 12'd4095;
            12'd2913: current_page <= 12'd4095;
            12'd2914: current_page <= 12'd4095;
            12'd2915: current_page <= 12'd4095;
            12'd2916: current_page <= 12'd4095;
            12'd2917: current_page <= 12'd4095;
            12'd2918: current_page <= 12'd4095;
            12'd2919: current_page <= 12'd4095;
            12'd2920: current_page <= 12'd4095;
            12'd2921: current_page <= 12'd4095;
            12'd2922: current_page <= 12'd4095;
            12'd2923: current_page <= 12'd4095;
            12'd2924: current_page <= 12'd4095;
            12'd2925: current_page <= 12'd4095;
            12'd2926: current_page <= 12'd4095;
            12'd2927: current_page <= 12'd4095;
            12'd2928: current_page <= 12'd4095;
            12'd2929: current_page <= 12'd4095;
            12'd2930: current_page <= 12'd4095;
            12'd2931: current_page <= 12'd4095;
            12'd2932: current_page <= 12'd4095;
            12'd2933: current_page <= 12'd4095;
            12'd2934: current_page <= 12'd4095;
            12'd2935: current_page <= 12'd4095;
            12'd2936: current_page <= 12'd4095;
            12'd2937: current_page <= 12'd4095;
            12'd2938: current_page <= 12'd4095;
            12'd2939: current_page <= 12'd4095;
            12'd2940: current_page <= 12'd4095;
            12'd2941: current_page <= 12'd4095;
            12'd2942: current_page <= 12'd4095;
            12'd2943: current_page <= 12'd4095;
            12'd2944: current_page <= 12'd4095;
            12'd2945: current_page <= 12'd4095;
            12'd2946: current_page <= 12'd4095;
            12'd2947: current_page <= 12'd4095;
            12'd2948: current_page <= 12'd4095;
            12'd2949: current_page <= 12'd4095;
            12'd2950: current_page <= 12'd4095;
            12'd2951: current_page <= 12'd4095;
            12'd2952: current_page <= 12'd4095;
            12'd2953: current_page <= 12'd4095;
            12'd2954: current_page <= 12'd4095;
            12'd2955: current_page <= 12'd4095;
            12'd2956: current_page <= 12'd4095;
            12'd2957: current_page <= 12'd4095;
            12'd2958: current_page <= 12'd4095;
            12'd2959: current_page <= 12'd4095;
            12'd2960: current_page <= 12'd4095;
            12'd2961: current_page <= 12'd4095;
            12'd2962: current_page <= 12'd4095;
            12'd2963: current_page <= 12'd4095;
            12'd2964: current_page <= 12'd4095;
            12'd2965: current_page <= 12'd4095;
            12'd2966: current_page <= 12'd4095;
            12'd2967: current_page <= 12'd4095;
            12'd2968: current_page <= 12'd4095;
            12'd2969: current_page <= 12'd4095;
            12'd2970: current_page <= 12'd4095;
            12'd2971: current_page <= 12'd4095;
            12'd2972: current_page <= 12'd4095;
            12'd2973: current_page <= 12'd4095;
            12'd2974: current_page <= 12'd4095;
            12'd2975: current_page <= 12'd4095;
            12'd2976: current_page <= 12'd4095;
            12'd2977: current_page <= 12'd4095;
            12'd2978: current_page <= 12'd4095;
            12'd2979: current_page <= 12'd4095;
            12'd2980: current_page <= 12'd4095;
            12'd2981: current_page <= 12'd4095;
            12'd2982: current_page <= 12'd4095;
            12'd2983: current_page <= 12'd4095;
            12'd2984: current_page <= 12'd4095;
            12'd2985: current_page <= 12'd4095;
            12'd2986: current_page <= 12'd4095;
            12'd2987: current_page <= 12'd4095;
            12'd2988: current_page <= 12'd4095;
            12'd2989: current_page <= 12'd4095;
            12'd2990: current_page <= 12'd4095;
            12'd2991: current_page <= 12'd4095;
            12'd2992: current_page <= 12'd4095;
            12'd2993: current_page <= 12'd4095;
            12'd2994: current_page <= 12'd4095;
            12'd2995: current_page <= 12'd4095;
            12'd2996: current_page <= 12'd4095;
            12'd2997: current_page <= 12'd4095;
            12'd2998: current_page <= 12'd4095;
            12'd2999: current_page <= 12'd4095;
            12'd3000: current_page <= 12'd4095;
            12'd3001: current_page <= 12'd4095;
            12'd3002: current_page <= 12'd4095;
            12'd3003: current_page <= 12'd4095;
            12'd3004: current_page <= 12'd4095;
            12'd3005: current_page <= 12'd4095;
            12'd3006: current_page <= 12'd4095;
            12'd3007: current_page <= 12'd4095;
            12'd3008: current_page <= 12'd4095;
            12'd3009: current_page <= 12'd4095;
            12'd3010: current_page <= 12'd4095;
            12'd3011: current_page <= 12'd4095;
            12'd3012: current_page <= 12'd4095;
            12'd3013: current_page <= 12'd4095;
            12'd3014: current_page <= 12'd4095;
            12'd3015: current_page <= 12'd4095;
            12'd3016: current_page <= 12'd4095;
            12'd3017: current_page <= 12'd4095;
            12'd3018: current_page <= 12'd4095;
            12'd3019: current_page <= 12'd4095;
            12'd3020: current_page <= 12'd4095;
            12'd3021: current_page <= 12'd4095;
            12'd3022: current_page <= 12'd4095;
            12'd3023: current_page <= 12'd4095;
            12'd3024: current_page <= 12'd4095;
            12'd3025: current_page <= 12'd4095;
            12'd3026: current_page <= 12'd4095;
            12'd3027: current_page <= 12'd4095;
            12'd3028: current_page <= 12'd4095;
            12'd3029: current_page <= 12'd4095;
            12'd3030: current_page <= 12'd4095;
            12'd3031: current_page <= 12'd4095;
            12'd3032: current_page <= 12'd4095;
            12'd3033: current_page <= 12'd4095;
            12'd3034: current_page <= 12'd4095;
            12'd3035: current_page <= 12'd4095;
            12'd3036: current_page <= 12'd4095;
            12'd3037: current_page <= 12'd4095;
            12'd3038: current_page <= 12'd4095;
            12'd3039: current_page <= 12'd4095;
            12'd3040: current_page <= 12'd4095;
            12'd3041: current_page <= 12'd4095;
            12'd3042: current_page <= 12'd4095;
            12'd3043: current_page <= 12'd4095;
            12'd3044: current_page <= 12'd4095;
            12'd3045: current_page <= 12'd4095;
            12'd3046: current_page <= 12'd4095;
            12'd3047: current_page <= 12'd4095;
            12'd3048: current_page <= 12'd4095;
            12'd3049: current_page <= 12'd4095;
            12'd3050: current_page <= 12'd4095;
            12'd3051: current_page <= 12'd4095;
            12'd3052: current_page <= 12'd4095;
            12'd3053: current_page <= 12'd4095;
            12'd3054: current_page <= 12'd4095;
            12'd3055: current_page <= 12'd4095;
            12'd3056: current_page <= 12'd4095;
            12'd3057: current_page <= 12'd4095;
            12'd3058: current_page <= 12'd4095;
            12'd3059: current_page <= 12'd4095;
            12'd3060: current_page <= 12'd4095;
            12'd3061: current_page <= 12'd4095;
            12'd3062: current_page <= 12'd4095;
            12'd3063: current_page <= 12'd4095;
            12'd3064: current_page <= 12'd4095;
            12'd3065: current_page <= 12'd4095;
            12'd3066: current_page <= 12'd4095;
            12'd3067: current_page <= 12'd4095;
            12'd3068: current_page <= 12'd4095;
            12'd3069: current_page <= 12'd4095;
            12'd3070: current_page <= 12'd4095;
            12'd3071: current_page <= 12'd4095;
            12'd3072: current_page <= 12'd4095;
            12'd3073: current_page <= 12'd4095;
            12'd3074: current_page <= 12'd4095;
            12'd3075: current_page <= 12'd4095;
            12'd3076: current_page <= 12'd4095;
            12'd3077: current_page <= 12'd4095;
            12'd3078: current_page <= 12'd4095;
            12'd3079: current_page <= 12'd4095;
            12'd3080: current_page <= 12'd4095;
            12'd3081: current_page <= 12'd4095;
            12'd3082: current_page <= 12'd4095;
            12'd3083: current_page <= 12'd4095;
            12'd3084: current_page <= 12'd4095;
            12'd3085: current_page <= 12'd4095;
            12'd3086: current_page <= 12'd4095;
            12'd3087: current_page <= 12'd4095;
            12'd3088: current_page <= 12'd4095;
            12'd3089: current_page <= 12'd4095;
            12'd3090: current_page <= 12'd4095;
            12'd3091: current_page <= 12'd4095;
            12'd3092: current_page <= 12'd4095;
            12'd3093: current_page <= 12'd4095;
            12'd3094: current_page <= 12'd4095;
            12'd3095: current_page <= 12'd4095;
            12'd3096: current_page <= 12'd4095;
            12'd3097: current_page <= 12'd4095;
            12'd3098: current_page <= 12'd4095;
            12'd3099: current_page <= 12'd4095;
            12'd3100: current_page <= 12'd4095;
            12'd3101: current_page <= 12'd4095;
            12'd3102: current_page <= 12'd4095;
            12'd3103: current_page <= 12'd4095;
            12'd3104: current_page <= 12'd4095;
            12'd3105: current_page <= 12'd4095;
            12'd3106: current_page <= 12'd4095;
            12'd3107: current_page <= 12'd4095;
            12'd3108: current_page <= 12'd4095;
            12'd3109: current_page <= 12'd4095;
            12'd3110: current_page <= 12'd4095;
            12'd3111: current_page <= 12'd4095;
            12'd3112: current_page <= 12'd4095;
            12'd3113: current_page <= 12'd4095;
            12'd3114: current_page <= 12'd4095;
            12'd3115: current_page <= 12'd4095;
            12'd3116: current_page <= 12'd4095;
            12'd3117: current_page <= 12'd4095;
            12'd3118: current_page <= 12'd4095;
            12'd3119: current_page <= 12'd4095;
            12'd3120: current_page <= 12'd4095;
            12'd3121: current_page <= 12'd4095;
            12'd3122: current_page <= 12'd4095;
            12'd3123: current_page <= 12'd4095;
            12'd3124: current_page <= 12'd4095;
            12'd3125: current_page <= 12'd4095;
            12'd3126: current_page <= 12'd4095;
            12'd3127: current_page <= 12'd4095;
            12'd3128: current_page <= 12'd4095;
            12'd3129: current_page <= 12'd4095;
            12'd3130: current_page <= 12'd4095;
            12'd3131: current_page <= 12'd4095;
            12'd3132: current_page <= 12'd4095;
            12'd3133: current_page <= 12'd4095;
            12'd3134: current_page <= 12'd4095;
            12'd3135: current_page <= 12'd4095;
            12'd3136: current_page <= 12'd4095;
            12'd3137: current_page <= 12'd4095;
            12'd3138: current_page <= 12'd4095;
            12'd3139: current_page <= 12'd4095;
            12'd3140: current_page <= 12'd4095;
            12'd3141: current_page <= 12'd4095;
            12'd3142: current_page <= 12'd4095;
            12'd3143: current_page <= 12'd4095;
            12'd3144: current_page <= 12'd4095;
            12'd3145: current_page <= 12'd4095;
            12'd3146: current_page <= 12'd4095;
            12'd3147: current_page <= 12'd4095;
            12'd3148: current_page <= 12'd4095;
            12'd3149: current_page <= 12'd4095;
            12'd3150: current_page <= 12'd4095;
            12'd3151: current_page <= 12'd4095;
            12'd3152: current_page <= 12'd4095;
            12'd3153: current_page <= 12'd4095;
            12'd3154: current_page <= 12'd4095;
            12'd3155: current_page <= 12'd4095;
            12'd3156: current_page <= 12'd4095;
            12'd3157: current_page <= 12'd4095;
            12'd3158: current_page <= 12'd4095;
            12'd3159: current_page <= 12'd4095;
            12'd3160: current_page <= 12'd4095;
            12'd3161: current_page <= 12'd4095;
            12'd3162: current_page <= 12'd4095;
            12'd3163: current_page <= 12'd4095;
            12'd3164: current_page <= 12'd4095;
            12'd3165: current_page <= 12'd4095;
            12'd3166: current_page <= 12'd4095;
            12'd3167: current_page <= 12'd4095;
            12'd3168: current_page <= 12'd4095;
            12'd3169: current_page <= 12'd4095;
            12'd3170: current_page <= 12'd4095;
            12'd3171: current_page <= 12'd4095;
            12'd3172: current_page <= 12'd4095;
            12'd3173: current_page <= 12'd4095;
            12'd3174: current_page <= 12'd4095;
            12'd3175: current_page <= 12'd4095;
            12'd3176: current_page <= 12'd4095;
            12'd3177: current_page <= 12'd4095;
            12'd3178: current_page <= 12'd4095;
            12'd3179: current_page <= 12'd4095;
            12'd3180: current_page <= 12'd4095;
            12'd3181: current_page <= 12'd4095;
            12'd3182: current_page <= 12'd4095;
            12'd3183: current_page <= 12'd4095;
            12'd3184: current_page <= 12'd4095;
            12'd3185: current_page <= 12'd4095;
            12'd3186: current_page <= 12'd4095;
            12'd3187: current_page <= 12'd4095;
            12'd3188: current_page <= 12'd4095;
            12'd3189: current_page <= 12'd4095;
            12'd3190: current_page <= 12'd4095;
            12'd3191: current_page <= 12'd4095;
            12'd3192: current_page <= 12'd4095;
            12'd3193: current_page <= 12'd4095;
            12'd3194: current_page <= 12'd4095;
            12'd3195: current_page <= 12'd4095;
            12'd3196: current_page <= 12'd4095;
            12'd3197: current_page <= 12'd4095;
            12'd3198: current_page <= 12'd4095;
            12'd3199: current_page <= 12'd4095;
            12'd3200: current_page <= 12'd4095;
            12'd3201: current_page <= 12'd4095;
            12'd3202: current_page <= 12'd4095;
            12'd3203: current_page <= 12'd4095;
            12'd3204: current_page <= 12'd4095;
            12'd3205: current_page <= 12'd4095;
            12'd3206: current_page <= 12'd4095;
            12'd3207: current_page <= 12'd4095;
            12'd3208: current_page <= 12'd4095;
            12'd3209: current_page <= 12'd4095;
            12'd3210: current_page <= 12'd4095;
            12'd3211: current_page <= 12'd4095;
            12'd3212: current_page <= 12'd4095;
            12'd3213: current_page <= 12'd4095;
            12'd3214: current_page <= 12'd4095;
            12'd3215: current_page <= 12'd4095;
            12'd3216: current_page <= 12'd4095;
            12'd3217: current_page <= 12'd4095;
            12'd3218: current_page <= 12'd4095;
            12'd3219: current_page <= 12'd4095;
            12'd3220: current_page <= 12'd4095;
            12'd3221: current_page <= 12'd4095;
            12'd3222: current_page <= 12'd4095;
            12'd3223: current_page <= 12'd4095;
            12'd3224: current_page <= 12'd4095;
            12'd3225: current_page <= 12'd4095;
            12'd3226: current_page <= 12'd4095;
            12'd3227: current_page <= 12'd4095;
            12'd3228: current_page <= 12'd4095;
            12'd3229: current_page <= 12'd4095;
            12'd3230: current_page <= 12'd4095;
            12'd3231: current_page <= 12'd4095;
            12'd3232: current_page <= 12'd4095;
            12'd3233: current_page <= 12'd4095;
            12'd3234: current_page <= 12'd4095;
            12'd3235: current_page <= 12'd4095;
            12'd3236: current_page <= 12'd4095;
            12'd3237: current_page <= 12'd4095;
            12'd3238: current_page <= 12'd4095;
            12'd3239: current_page <= 12'd4095;
            12'd3240: current_page <= 12'd4095;
            12'd3241: current_page <= 12'd4095;
            12'd3242: current_page <= 12'd4095;
            12'd3243: current_page <= 12'd4095;
            12'd3244: current_page <= 12'd4095;
            12'd3245: current_page <= 12'd4095;
            12'd3246: current_page <= 12'd4095;
            12'd3247: current_page <= 12'd4095;
            12'd3248: current_page <= 12'd4095;
            12'd3249: current_page <= 12'd4095;
            12'd3250: current_page <= 12'd4095;
            12'd3251: current_page <= 12'd4095;
            12'd3252: current_page <= 12'd4095;
            12'd3253: current_page <= 12'd4095;
            12'd3254: current_page <= 12'd4095;
            12'd3255: current_page <= 12'd4095;
            12'd3256: current_page <= 12'd4095;
            12'd3257: current_page <= 12'd4095;
            12'd3258: current_page <= 12'd4095;
            12'd3259: current_page <= 12'd4095;
            12'd3260: current_page <= 12'd4095;
            12'd3261: current_page <= 12'd4095;
            12'd3262: current_page <= 12'd4095;
            12'd3263: current_page <= 12'd4095;
            12'd3264: current_page <= 12'd4095;
            12'd3265: current_page <= 12'd4095;
            12'd3266: current_page <= 12'd4095;
            12'd3267: current_page <= 12'd4095;
            12'd3268: current_page <= 12'd4095;
            12'd3269: current_page <= 12'd4095;
            12'd3270: current_page <= 12'd4095;
            12'd3271: current_page <= 12'd4095;
            12'd3272: current_page <= 12'd4095;
            12'd3273: current_page <= 12'd4095;
            12'd3274: current_page <= 12'd4095;
            12'd3275: current_page <= 12'd4095;
            12'd3276: current_page <= 12'd4095;
            12'd3277: current_page <= 12'd4095;
            12'd3278: current_page <= 12'd4095;
            12'd3279: current_page <= 12'd4095;
            12'd3280: current_page <= 12'd4095;
            12'd3281: current_page <= 12'd4095;
            12'd3282: current_page <= 12'd4095;
            12'd3283: current_page <= 12'd4095;
            12'd3284: current_page <= 12'd4095;
            12'd3285: current_page <= 12'd4095;
            12'd3286: current_page <= 12'd4095;
            12'd3287: current_page <= 12'd4095;
            12'd3288: current_page <= 12'd4095;
            12'd3289: current_page <= 12'd4095;
            12'd3290: current_page <= 12'd4095;
            12'd3291: current_page <= 12'd4095;
            12'd3292: current_page <= 12'd4095;
            12'd3293: current_page <= 12'd4095;
            12'd3294: current_page <= 12'd4095;
            12'd3295: current_page <= 12'd4095;
            12'd3296: current_page <= 12'd4095;
            12'd3297: current_page <= 12'd4095;
            12'd3298: current_page <= 12'd4095;
            12'd3299: current_page <= 12'd4095;
            12'd3300: current_page <= 12'd4095;
            12'd3301: current_page <= 12'd4095;
            12'd3302: current_page <= 12'd4095;
            12'd3303: current_page <= 12'd4095;
            12'd3304: current_page <= 12'd4095;
            12'd3305: current_page <= 12'd4095;
            12'd3306: current_page <= 12'd4095;
            12'd3307: current_page <= 12'd4095;
            12'd3308: current_page <= 12'd4095;
            12'd3309: current_page <= 12'd4095;
            12'd3310: current_page <= 12'd4095;
            12'd3311: current_page <= 12'd4095;
            12'd3312: current_page <= 12'd4095;
            12'd3313: current_page <= 12'd4095;
            12'd3314: current_page <= 12'd4095;
            12'd3315: current_page <= 12'd4095;
            12'd3316: current_page <= 12'd4095;
            12'd3317: current_page <= 12'd4095;
            12'd3318: current_page <= 12'd4095;
            12'd3319: current_page <= 12'd4095;
            12'd3320: current_page <= 12'd4095;
            12'd3321: current_page <= 12'd4095;
            12'd3322: current_page <= 12'd4095;
            12'd3323: current_page <= 12'd4095;
            12'd3324: current_page <= 12'd4095;
            12'd3325: current_page <= 12'd4095;
            12'd3326: current_page <= 12'd4095;
            12'd3327: current_page <= 12'd4095;
            12'd3328: current_page <= 12'd4095;
            12'd3329: current_page <= 12'd4095;
            12'd3330: current_page <= 12'd4095;
            12'd3331: current_page <= 12'd4095;
            12'd3332: current_page <= 12'd4095;
            12'd3333: current_page <= 12'd4095;
            12'd3334: current_page <= 12'd4095;
            12'd3335: current_page <= 12'd4095;
            12'd3336: current_page <= 12'd4095;
            12'd3337: current_page <= 12'd4095;
            12'd3338: current_page <= 12'd4095;
            12'd3339: current_page <= 12'd4095;
            12'd3340: current_page <= 12'd4095;
            12'd3341: current_page <= 12'd4095;
            12'd3342: current_page <= 12'd4095;
            12'd3343: current_page <= 12'd4095;
            12'd3344: current_page <= 12'd4095;
            12'd3345: current_page <= 12'd4095;
            12'd3346: current_page <= 12'd4095;
            12'd3347: current_page <= 12'd4095;
            12'd3348: current_page <= 12'd4095;
            12'd3349: current_page <= 12'd4095;
            12'd3350: current_page <= 12'd4095;
            12'd3351: current_page <= 12'd4095;
            12'd3352: current_page <= 12'd4095;
            12'd3353: current_page <= 12'd4095;
            12'd3354: current_page <= 12'd4095;
            12'd3355: current_page <= 12'd4095;
            12'd3356: current_page <= 12'd4095;
            12'd3357: current_page <= 12'd4095;
            12'd3358: current_page <= 12'd4095;
            12'd3359: current_page <= 12'd4095;
            12'd3360: current_page <= 12'd4095;
            12'd3361: current_page <= 12'd4095;
            12'd3362: current_page <= 12'd4095;
            12'd3363: current_page <= 12'd4095;
            12'd3364: current_page <= 12'd4095;
            12'd3365: current_page <= 12'd4095;
            12'd3366: current_page <= 12'd4095;
            12'd3367: current_page <= 12'd4095;
            12'd3368: current_page <= 12'd4095;
            12'd3369: current_page <= 12'd4095;
            12'd3370: current_page <= 12'd4095;
            12'd3371: current_page <= 12'd4095;
            12'd3372: current_page <= 12'd4095;
            12'd3373: current_page <= 12'd4095;
            12'd3374: current_page <= 12'd4095;
            12'd3375: current_page <= 12'd4095;
            12'd3376: current_page <= 12'd4095;
            12'd3377: current_page <= 12'd4095;
            12'd3378: current_page <= 12'd4095;
            12'd3379: current_page <= 12'd4095;
            12'd3380: current_page <= 12'd4095;
            12'd3381: current_page <= 12'd4095;
            12'd3382: current_page <= 12'd4095;
            12'd3383: current_page <= 12'd4095;
            12'd3384: current_page <= 12'd4095;
            12'd3385: current_page <= 12'd4095;
            12'd3386: current_page <= 12'd4095;
            12'd3387: current_page <= 12'd4095;
            12'd3388: current_page <= 12'd4095;
            12'd3389: current_page <= 12'd4095;
            12'd3390: current_page <= 12'd4095;
            12'd3391: current_page <= 12'd4095;
            12'd3392: current_page <= 12'd4095;
            12'd3393: current_page <= 12'd4095;
            12'd3394: current_page <= 12'd4095;
            12'd3395: current_page <= 12'd4095;
            12'd3396: current_page <= 12'd4095;
            12'd3397: current_page <= 12'd4095;
            12'd3398: current_page <= 12'd4095;
            12'd3399: current_page <= 12'd4095;
            12'd3400: current_page <= 12'd4095;
            12'd3401: current_page <= 12'd4095;
            12'd3402: current_page <= 12'd4095;
            12'd3403: current_page <= 12'd4095;
            12'd3404: current_page <= 12'd4095;
            12'd3405: current_page <= 12'd4095;
            12'd3406: current_page <= 12'd4095;
            12'd3407: current_page <= 12'd4095;
            12'd3408: current_page <= 12'd4095;
            12'd3409: current_page <= 12'd4095;
            12'd3410: current_page <= 12'd4095;
            12'd3411: current_page <= 12'd4095;
            12'd3412: current_page <= 12'd4095;
            12'd3413: current_page <= 12'd4095;
            12'd3414: current_page <= 12'd4095;
            12'd3415: current_page <= 12'd4095;
            12'd3416: current_page <= 12'd4095;
            12'd3417: current_page <= 12'd4095;
            12'd3418: current_page <= 12'd4095;
            12'd3419: current_page <= 12'd4095;
            12'd3420: current_page <= 12'd4095;
            12'd3421: current_page <= 12'd4095;
            12'd3422: current_page <= 12'd4095;
            12'd3423: current_page <= 12'd4095;
            12'd3424: current_page <= 12'd4095;
            12'd3425: current_page <= 12'd4095;
            12'd3426: current_page <= 12'd4095;
            12'd3427: current_page <= 12'd4095;
            12'd3428: current_page <= 12'd4095;
            12'd3429: current_page <= 12'd4095;
            12'd3430: current_page <= 12'd4095;
            12'd3431: current_page <= 12'd4095;
            12'd3432: current_page <= 12'd4095;
            12'd3433: current_page <= 12'd4095;
            12'd3434: current_page <= 12'd4095;
            12'd3435: current_page <= 12'd4095;
            12'd3436: current_page <= 12'd4095;
            12'd3437: current_page <= 12'd4095;
            12'd3438: current_page <= 12'd4095;
            12'd3439: current_page <= 12'd4095;
            12'd3440: current_page <= 12'd4095;
            12'd3441: current_page <= 12'd4095;
            12'd3442: current_page <= 12'd4095;
            12'd3443: current_page <= 12'd4095;
            12'd3444: current_page <= 12'd4095;
            12'd3445: current_page <= 12'd4095;
            12'd3446: current_page <= 12'd4095;
            12'd3447: current_page <= 12'd4095;
            12'd3448: current_page <= 12'd4095;
            12'd3449: current_page <= 12'd4095;
            12'd3450: current_page <= 12'd4095;
            12'd3451: current_page <= 12'd4095;
            12'd3452: current_page <= 12'd4095;
            12'd3453: current_page <= 12'd4095;
            12'd3454: current_page <= 12'd4095;
            12'd3455: current_page <= 12'd4095;
            12'd3456: current_page <= 12'd4095;
            12'd3457: current_page <= 12'd4095;
            12'd3458: current_page <= 12'd4095;
            12'd3459: current_page <= 12'd4095;
            12'd3460: current_page <= 12'd4095;
            12'd3461: current_page <= 12'd4095;
            12'd3462: current_page <= 12'd4095;
            12'd3463: current_page <= 12'd4095;
            12'd3464: current_page <= 12'd4095;
            12'd3465: current_page <= 12'd4095;
            12'd3466: current_page <= 12'd4095;
            12'd3467: current_page <= 12'd4095;
            12'd3468: current_page <= 12'd4095;
            12'd3469: current_page <= 12'd4095;
            12'd3470: current_page <= 12'd4095;
            12'd3471: current_page <= 12'd4095;
            12'd3472: current_page <= 12'd4095;
            12'd3473: current_page <= 12'd4095;
            12'd3474: current_page <= 12'd4095;
            12'd3475: current_page <= 12'd4095;
            12'd3476: current_page <= 12'd4095;
            12'd3477: current_page <= 12'd4095;
            12'd3478: current_page <= 12'd4095;
            12'd3479: current_page <= 12'd4095;
            12'd3480: current_page <= 12'd4095;
            12'd3481: current_page <= 12'd4095;
            12'd3482: current_page <= 12'd4095;
            12'd3483: current_page <= 12'd4095;
            12'd3484: current_page <= 12'd4095;
            12'd3485: current_page <= 12'd4095;
            12'd3486: current_page <= 12'd4095;
            12'd3487: current_page <= 12'd4095;
            12'd3488: current_page <= 12'd4095;
            12'd3489: current_page <= 12'd4095;
            12'd3490: current_page <= 12'd4095;
            12'd3491: current_page <= 12'd4095;
            12'd3492: current_page <= 12'd4095;
            12'd3493: current_page <= 12'd4095;
            12'd3494: current_page <= 12'd4095;
            12'd3495: current_page <= 12'd4095;
            12'd3496: current_page <= 12'd4095;
            12'd3497: current_page <= 12'd4095;
            12'd3498: current_page <= 12'd4095;
            12'd3499: current_page <= 12'd4095;
            12'd3500: current_page <= 12'd4095;
            12'd3501: current_page <= 12'd4095;
            12'd3502: current_page <= 12'd4095;
            12'd3503: current_page <= 12'd4095;
            12'd3504: current_page <= 12'd4095;
            12'd3505: current_page <= 12'd4095;
            12'd3506: current_page <= 12'd4095;
            12'd3507: current_page <= 12'd4095;
            12'd3508: current_page <= 12'd4095;
            12'd3509: current_page <= 12'd4095;
            12'd3510: current_page <= 12'd4095;
            12'd3511: current_page <= 12'd4095;
            12'd3512: current_page <= 12'd4095;
            12'd3513: current_page <= 12'd4095;
            12'd3514: current_page <= 12'd4095;
            12'd3515: current_page <= 12'd4095;
            12'd3516: current_page <= 12'd4095;
            12'd3517: current_page <= 12'd4095;
            12'd3518: current_page <= 12'd4095;
            12'd3519: current_page <= 12'd4095;
            12'd3520: current_page <= 12'd4095;
            12'd3521: current_page <= 12'd4095;
            12'd3522: current_page <= 12'd4095;
            12'd3523: current_page <= 12'd4095;
            12'd3524: current_page <= 12'd4095;
            12'd3525: current_page <= 12'd4095;
            12'd3526: current_page <= 12'd4095;
            12'd3527: current_page <= 12'd4095;
            12'd3528: current_page <= 12'd4095;
            12'd3529: current_page <= 12'd4095;
            12'd3530: current_page <= 12'd4095;
            12'd3531: current_page <= 12'd4095;
            12'd3532: current_page <= 12'd4095;
            12'd3533: current_page <= 12'd4095;
            12'd3534: current_page <= 12'd4095;
            12'd3535: current_page <= 12'd4095;
            12'd3536: current_page <= 12'd4095;
            12'd3537: current_page <= 12'd4095;
            12'd3538: current_page <= 12'd4095;
            12'd3539: current_page <= 12'd4095;
            12'd3540: current_page <= 12'd4095;
            12'd3541: current_page <= 12'd4095;
            12'd3542: current_page <= 12'd4095;
            12'd3543: current_page <= 12'd4095;
            12'd3544: current_page <= 12'd4095;
            12'd3545: current_page <= 12'd4095;
            12'd3546: current_page <= 12'd4095;
            12'd3547: current_page <= 12'd4095;
            12'd3548: current_page <= 12'd4095;
            12'd3549: current_page <= 12'd4095;
            12'd3550: current_page <= 12'd4095;
            12'd3551: current_page <= 12'd4095;
            12'd3552: current_page <= 12'd4095;
            12'd3553: current_page <= 12'd4095;
            12'd3554: current_page <= 12'd4095;
            12'd3555: current_page <= 12'd4095;
            12'd3556: current_page <= 12'd4095;
            12'd3557: current_page <= 12'd4095;
            12'd3558: current_page <= 12'd4095;
            12'd3559: current_page <= 12'd4095;
            12'd3560: current_page <= 12'd4095;
            12'd3561: current_page <= 12'd4095;
            12'd3562: current_page <= 12'd4095;
            12'd3563: current_page <= 12'd4095;
            12'd3564: current_page <= 12'd4095;
            12'd3565: current_page <= 12'd4095;
            12'd3566: current_page <= 12'd4095;
            12'd3567: current_page <= 12'd4095;
            12'd3568: current_page <= 12'd4095;
            12'd3569: current_page <= 12'd4095;
            12'd3570: current_page <= 12'd4095;
            12'd3571: current_page <= 12'd4095;
            12'd3572: current_page <= 12'd4095;
            12'd3573: current_page <= 12'd4095;
            12'd3574: current_page <= 12'd4095;
            12'd3575: current_page <= 12'd4095;
            12'd3576: current_page <= 12'd4095;
            12'd3577: current_page <= 12'd4095;
            12'd3578: current_page <= 12'd4095;
            12'd3579: current_page <= 12'd4095;
            12'd3580: current_page <= 12'd4095;
            12'd3581: current_page <= 12'd4095;
            12'd3582: current_page <= 12'd4095;
            12'd3583: current_page <= 12'd4095;
            12'd3584: current_page <= 12'd4095;
            12'd3585: current_page <= 12'd4095;
            12'd3586: current_page <= 12'd4095;
            12'd3587: current_page <= 12'd4095;
            12'd3588: current_page <= 12'd4095;
            12'd3589: current_page <= 12'd4095;
            12'd3590: current_page <= 12'd4095;
            12'd3591: current_page <= 12'd4095;
            12'd3592: current_page <= 12'd4095;
            12'd3593: current_page <= 12'd4095;
            12'd3594: current_page <= 12'd4095;
            12'd3595: current_page <= 12'd4095;
            12'd3596: current_page <= 12'd4095;
            12'd3597: current_page <= 12'd4095;
            12'd3598: current_page <= 12'd4095;
            12'd3599: current_page <= 12'd4095;
            12'd3600: current_page <= 12'd4095;
            12'd3601: current_page <= 12'd4095;
            12'd3602: current_page <= 12'd4095;
            12'd3603: current_page <= 12'd4095;
            12'd3604: current_page <= 12'd4095;
            12'd3605: current_page <= 12'd4095;
            12'd3606: current_page <= 12'd4095;
            12'd3607: current_page <= 12'd4095;
            12'd3608: current_page <= 12'd4095;
            12'd3609: current_page <= 12'd4095;
            12'd3610: current_page <= 12'd4095;
            12'd3611: current_page <= 12'd4095;
            12'd3612: current_page <= 12'd4095;
            12'd3613: current_page <= 12'd4095;
            12'd3614: current_page <= 12'd4095;
            12'd3615: current_page <= 12'd4095;
            12'd3616: current_page <= 12'd4095;
            12'd3617: current_page <= 12'd4095;
            12'd3618: current_page <= 12'd4095;
            12'd3619: current_page <= 12'd4095;
            12'd3620: current_page <= 12'd4095;
            12'd3621: current_page <= 12'd4095;
            12'd3622: current_page <= 12'd4095;
            12'd3623: current_page <= 12'd4095;
            12'd3624: current_page <= 12'd4095;
            12'd3625: current_page <= 12'd4095;
            12'd3626: current_page <= 12'd4095;
            12'd3627: current_page <= 12'd4095;
            12'd3628: current_page <= 12'd4095;
            12'd3629: current_page <= 12'd4095;
            12'd3630: current_page <= 12'd4095;
            12'd3631: current_page <= 12'd4095;
            12'd3632: current_page <= 12'd4095;
            12'd3633: current_page <= 12'd4095;
            12'd3634: current_page <= 12'd4095;
            12'd3635: current_page <= 12'd4095;
            12'd3636: current_page <= 12'd4095;
            12'd3637: current_page <= 12'd4095;
            12'd3638: current_page <= 12'd4095;
            12'd3639: current_page <= 12'd4095;
            12'd3640: current_page <= 12'd4095;
            12'd3641: current_page <= 12'd4095;
            12'd3642: current_page <= 12'd4095;
            12'd3643: current_page <= 12'd4095;
            12'd3644: current_page <= 12'd4095;
            12'd3645: current_page <= 12'd4095;
            12'd3646: current_page <= 12'd4095;
            12'd3647: current_page <= 12'd4095;
            12'd3648: current_page <= 12'd4095;
            12'd3649: current_page <= 12'd4095;
            12'd3650: current_page <= 12'd4095;
            12'd3651: current_page <= 12'd4095;
            12'd3652: current_page <= 12'd4095;
            12'd3653: current_page <= 12'd4095;
            12'd3654: current_page <= 12'd4095;
            12'd3655: current_page <= 12'd4095;
            12'd3656: current_page <= 12'd4095;
            12'd3657: current_page <= 12'd4095;
            12'd3658: current_page <= 12'd4095;
            12'd3659: current_page <= 12'd4095;
            12'd3660: current_page <= 12'd4095;
            12'd3661: current_page <= 12'd4095;
            12'd3662: current_page <= 12'd4095;
            12'd3663: current_page <= 12'd4095;
            12'd3664: current_page <= 12'd4095;
            12'd3665: current_page <= 12'd4095;
            12'd3666: current_page <= 12'd4095;
            12'd3667: current_page <= 12'd4095;
            12'd3668: current_page <= 12'd4095;
            12'd3669: current_page <= 12'd4095;
            12'd3670: current_page <= 12'd4095;
            12'd3671: current_page <= 12'd4095;
            12'd3672: current_page <= 12'd4095;
            12'd3673: current_page <= 12'd4095;
            12'd3674: current_page <= 12'd4095;
            12'd3675: current_page <= 12'd4095;
            12'd3676: current_page <= 12'd4095;
            12'd3677: current_page <= 12'd4095;
            12'd3678: current_page <= 12'd4095;
            12'd3679: current_page <= 12'd4095;
            12'd3680: current_page <= 12'd4095;
            12'd3681: current_page <= 12'd4095;
            12'd3682: current_page <= 12'd4095;
            12'd3683: current_page <= 12'd4095;
            12'd3684: current_page <= 12'd4095;
            12'd3685: current_page <= 12'd4095;
            12'd3686: current_page <= 12'd4095;
            12'd3687: current_page <= 12'd4095;
            12'd3688: current_page <= 12'd4095;
            12'd3689: current_page <= 12'd4095;
            12'd3690: current_page <= 12'd4095;
            12'd3691: current_page <= 12'd4095;
            12'd3692: current_page <= 12'd4095;
            12'd3693: current_page <= 12'd4095;
            12'd3694: current_page <= 12'd4095;
            12'd3695: current_page <= 12'd4095;
            12'd3696: current_page <= 12'd4095;
            12'd3697: current_page <= 12'd4095;
            12'd3698: current_page <= 12'd4095;
            12'd3699: current_page <= 12'd4095;
            12'd3700: current_page <= 12'd4095;
            12'd3701: current_page <= 12'd4095;
            12'd3702: current_page <= 12'd4095;
            12'd3703: current_page <= 12'd4095;
            12'd3704: current_page <= 12'd4095;
            12'd3705: current_page <= 12'd4095;
            12'd3706: current_page <= 12'd4095;
            12'd3707: current_page <= 12'd4095;
            12'd3708: current_page <= 12'd4095;
            12'd3709: current_page <= 12'd4095;
            12'd3710: current_page <= 12'd4095;
            12'd3711: current_page <= 12'd4095;
            12'd3712: current_page <= 12'd4095;
            12'd3713: current_page <= 12'd4095;
            12'd3714: current_page <= 12'd4095;
            12'd3715: current_page <= 12'd4095;
            12'd3716: current_page <= 12'd4095;
            12'd3717: current_page <= 12'd4095;
            12'd3718: current_page <= 12'd4095;
            12'd3719: current_page <= 12'd4095;
            12'd3720: current_page <= 12'd4095;
            12'd3721: current_page <= 12'd4095;
            12'd3722: current_page <= 12'd4095;
            12'd3723: current_page <= 12'd4095;
            12'd3724: current_page <= 12'd4095;
            12'd3725: current_page <= 12'd4095;
            12'd3726: current_page <= 12'd4095;
            12'd3727: current_page <= 12'd4095;
            12'd3728: current_page <= 12'd4095;
            12'd3729: current_page <= 12'd4095;
            12'd3730: current_page <= 12'd4095;
            12'd3731: current_page <= 12'd4095;
            12'd3732: current_page <= 12'd4095;
            12'd3733: current_page <= 12'd4095;
            12'd3734: current_page <= 12'd4095;
            12'd3735: current_page <= 12'd4095;
            12'd3736: current_page <= 12'd4095;
            12'd3737: current_page <= 12'd4095;
            12'd3738: current_page <= 12'd4095;
            12'd3739: current_page <= 12'd4095;
            12'd3740: current_page <= 12'd4095;
            12'd3741: current_page <= 12'd4095;
            12'd3742: current_page <= 12'd4095;
            12'd3743: current_page <= 12'd4095;
            12'd3744: current_page <= 12'd4095;
            12'd3745: current_page <= 12'd4095;
            12'd3746: current_page <= 12'd4095;
            12'd3747: current_page <= 12'd4095;
            12'd3748: current_page <= 12'd4095;
            12'd3749: current_page <= 12'd4095;
            12'd3750: current_page <= 12'd4095;
            12'd3751: current_page <= 12'd4095;
            12'd3752: current_page <= 12'd4095;
            12'd3753: current_page <= 12'd4095;
            12'd3754: current_page <= 12'd4095;
            12'd3755: current_page <= 12'd4095;
            12'd3756: current_page <= 12'd4095;
            12'd3757: current_page <= 12'd4095;
            12'd3758: current_page <= 12'd4095;
            12'd3759: current_page <= 12'd4095;
            12'd3760: current_page <= 12'd4095;
            12'd3761: current_page <= 12'd4095;
            12'd3762: current_page <= 12'd4095;
            12'd3763: current_page <= 12'd4095;
            12'd3764: current_page <= 12'd4095;
            12'd3765: current_page <= 12'd4095;
            12'd3766: current_page <= 12'd4095;
            12'd3767: current_page <= 12'd4095;
            12'd3768: current_page <= 12'd4095;
            12'd3769: current_page <= 12'd4095;
            12'd3770: current_page <= 12'd4095;
            12'd3771: current_page <= 12'd4095;
            12'd3772: current_page <= 12'd4095;
            12'd3773: current_page <= 12'd4095;
            12'd3774: current_page <= 12'd4095;
            12'd3775: current_page <= 12'd4095;
            12'd3776: current_page <= 12'd4095;
            12'd3777: current_page <= 12'd4095;
            12'd3778: current_page <= 12'd4095;
            12'd3779: current_page <= 12'd4095;
            12'd3780: current_page <= 12'd4095;
            12'd3781: current_page <= 12'd4095;
            12'd3782: current_page <= 12'd4095;
            12'd3783: current_page <= 12'd4095;
            12'd3784: current_page <= 12'd4095;
            12'd3785: current_page <= 12'd4095;
            12'd3786: current_page <= 12'd4095;
            12'd3787: current_page <= 12'd4095;
            12'd3788: current_page <= 12'd4095;
            12'd3789: current_page <= 12'd4095;
            12'd3790: current_page <= 12'd4095;
            12'd3791: current_page <= 12'd4095;
            12'd3792: current_page <= 12'd4095;
            12'd3793: current_page <= 12'd4095;
            12'd3794: current_page <= 12'd4095;
            12'd3795: current_page <= 12'd4095;
            12'd3796: current_page <= 12'd4095;
            12'd3797: current_page <= 12'd4095;
            12'd3798: current_page <= 12'd4095;
            12'd3799: current_page <= 12'd4095;
            12'd3800: current_page <= 12'd4095;
            12'd3801: current_page <= 12'd4095;
            12'd3802: current_page <= 12'd4095;
            12'd3803: current_page <= 12'd4095;
            12'd3804: current_page <= 12'd4095;
            12'd3805: current_page <= 12'd4095;
            12'd3806: current_page <= 12'd4095;
            12'd3807: current_page <= 12'd4095;
            12'd3808: current_page <= 12'd4095;
            12'd3809: current_page <= 12'd4095;
            12'd3810: current_page <= 12'd4095;
            12'd3811: current_page <= 12'd4095;
            12'd3812: current_page <= 12'd4095;
            12'd3813: current_page <= 12'd4095;
            12'd3814: current_page <= 12'd4095;
            12'd3815: current_page <= 12'd4095;
            12'd3816: current_page <= 12'd4095;
            12'd3817: current_page <= 12'd4095;
            12'd3818: current_page <= 12'd4095;
            12'd3819: current_page <= 12'd4095;
            12'd3820: current_page <= 12'd4095;
            12'd3821: current_page <= 12'd4095;
            12'd3822: current_page <= 12'd4095;
            12'd3823: current_page <= 12'd4095;
            12'd3824: current_page <= 12'd4095;
            12'd3825: current_page <= 12'd4095;
            12'd3826: current_page <= 12'd4095;
            12'd3827: current_page <= 12'd4095;
            12'd3828: current_page <= 12'd4095;
            12'd3829: current_page <= 12'd4095;
            12'd3830: current_page <= 12'd4095;
            12'd3831: current_page <= 12'd4095;
            12'd3832: current_page <= 12'd4095;
            12'd3833: current_page <= 12'd4095;
            12'd3834: current_page <= 12'd4095;
            12'd3835: current_page <= 12'd4095;
            12'd3836: current_page <= 12'd4095;
            12'd3837: current_page <= 12'd4095;
            12'd3838: current_page <= 12'd4095;
            12'd3839: current_page <= 12'd4095;
            12'd3840: current_page <= 12'd4095;
            12'd3841: current_page <= 12'd4095;
            12'd3842: current_page <= 12'd4095;
            12'd3843: current_page <= 12'd4095;
            12'd3844: current_page <= 12'd4095;
            12'd3845: current_page <= 12'd4095;
            12'd3846: current_page <= 12'd4095;
            12'd3847: current_page <= 12'd4095;
            12'd3848: current_page <= 12'd4095;
            12'd3849: current_page <= 12'd4095;
            12'd3850: current_page <= 12'd4095;
            12'd3851: current_page <= 12'd4095;
            12'd3852: current_page <= 12'd4095;
            12'd3853: current_page <= 12'd4095;
            12'd3854: current_page <= 12'd4095;
            12'd3855: current_page <= 12'd4095;
            12'd3856: current_page <= 12'd4095;
            12'd3857: current_page <= 12'd4095;
            12'd3858: current_page <= 12'd4095;
            12'd3859: current_page <= 12'd4095;
            12'd3860: current_page <= 12'd4095;
            12'd3861: current_page <= 12'd4095;
            12'd3862: current_page <= 12'd4095;
            12'd3863: current_page <= 12'd4095;
            12'd3864: current_page <= 12'd4095;
            12'd3865: current_page <= 12'd4095;
            12'd3866: current_page <= 12'd4095;
            12'd3867: current_page <= 12'd4095;
            12'd3868: current_page <= 12'd4095;
            12'd3869: current_page <= 12'd4095;
            12'd3870: current_page <= 12'd4095;
            12'd3871: current_page <= 12'd4095;
            12'd3872: current_page <= 12'd4095;
            12'd3873: current_page <= 12'd4095;
            12'd3874: current_page <= 12'd4095;
            12'd3875: current_page <= 12'd4095;
            12'd3876: current_page <= 12'd4095;
            12'd3877: current_page <= 12'd4095;
            12'd3878: current_page <= 12'd4095;
            12'd3879: current_page <= 12'd4095;
            12'd3880: current_page <= 12'd4095;
            12'd3881: current_page <= 12'd4095;
            12'd3882: current_page <= 12'd4095;
            12'd3883: current_page <= 12'd4095;
            12'd3884: current_page <= 12'd4095;
            12'd3885: current_page <= 12'd4095;
            12'd3886: current_page <= 12'd4095;
            12'd3887: current_page <= 12'd4095;
            12'd3888: current_page <= 12'd4095;
            12'd3889: current_page <= 12'd4095;
            12'd3890: current_page <= 12'd4095;
            12'd3891: current_page <= 12'd4095;
            12'd3892: current_page <= 12'd4095;
            12'd3893: current_page <= 12'd4095;
            12'd3894: current_page <= 12'd4095;
            12'd3895: current_page <= 12'd4095;
            12'd3896: current_page <= 12'd4095;
            12'd3897: current_page <= 12'd4095;
            12'd3898: current_page <= 12'd4095;
            12'd3899: current_page <= 12'd4095;
            12'd3900: current_page <= 12'd4095;
            12'd3901: current_page <= 12'd4095;
            12'd3902: current_page <= 12'd4095;
            12'd3903: current_page <= 12'd4095;
            12'd3904: current_page <= 12'd4095;
            12'd3905: current_page <= 12'd4095;
            12'd3906: current_page <= 12'd4095;
            12'd3907: current_page <= 12'd4095;
            12'd3908: current_page <= 12'd4095;
            12'd3909: current_page <= 12'd4095;
            12'd3910: current_page <= 12'd4095;
            12'd3911: current_page <= 12'd4095;
            12'd3912: current_page <= 12'd4095;
            12'd3913: current_page <= 12'd4095;
            12'd3914: current_page <= 12'd4095;
            12'd3915: current_page <= 12'd4095;
            12'd3916: current_page <= 12'd4095;
            12'd3917: current_page <= 12'd4095;
            12'd3918: current_page <= 12'd4095;
            12'd3919: current_page <= 12'd4095;
            12'd3920: current_page <= 12'd4095;
            12'd3921: current_page <= 12'd4095;
            12'd3922: current_page <= 12'd4095;
            12'd3923: current_page <= 12'd4095;
            12'd3924: current_page <= 12'd4095;
            12'd3925: current_page <= 12'd4095;
            12'd3926: current_page <= 12'd4095;
            12'd3927: current_page <= 12'd4095;
            12'd3928: current_page <= 12'd4095;
            12'd3929: current_page <= 12'd4095;
            12'd3930: current_page <= 12'd4095;
            12'd3931: current_page <= 12'd4095;
            12'd3932: current_page <= 12'd4095;
            12'd3933: current_page <= 12'd4095;
            12'd3934: current_page <= 12'd4095;
            12'd3935: current_page <= 12'd4095;
            12'd3936: current_page <= 12'd4095;
            12'd3937: current_page <= 12'd4095;
            12'd3938: current_page <= 12'd4095;
            12'd3939: current_page <= 12'd4095;
            12'd3940: current_page <= 12'd4095;
            12'd3941: current_page <= 12'd4095;
            12'd3942: current_page <= 12'd4095;
            12'd3943: current_page <= 12'd4095;
            12'd3944: current_page <= 12'd4095;
            12'd3945: current_page <= 12'd4095;
            12'd3946: current_page <= 12'd4095;
            12'd3947: current_page <= 12'd4095;
            12'd3948: current_page <= 12'd4095;
            12'd3949: current_page <= 12'd4095;
            12'd3950: current_page <= 12'd4095;
            12'd3951: current_page <= 12'd4095;
            12'd3952: current_page <= 12'd4095;
            12'd3953: current_page <= 12'd4095;
            12'd3954: current_page <= 12'd4095;
            12'd3955: current_page <= 12'd4095;
            12'd3956: current_page <= 12'd4095;
            12'd3957: current_page <= 12'd4095;
            12'd3958: current_page <= 12'd4095;
            12'd3959: current_page <= 12'd4095;
            12'd3960: current_page <= 12'd4095;
            12'd3961: current_page <= 12'd4095;
            12'd3962: current_page <= 12'd4095;
            12'd3963: current_page <= 12'd4095;
            12'd3964: current_page <= 12'd4095;
            12'd3965: current_page <= 12'd4095;
            12'd3966: current_page <= 12'd4095;
            12'd3967: current_page <= 12'd4095;
            12'd3968: current_page <= 12'd4095;
            12'd3969: current_page <= 12'd4095;
            12'd3970: current_page <= 12'd4095;
            12'd3971: current_page <= 12'd4095;
            12'd3972: current_page <= 12'd4095;
            12'd3973: current_page <= 12'd4095;
            12'd3974: current_page <= 12'd4095;
            12'd3975: current_page <= 12'd4095;
            12'd3976: current_page <= 12'd4095;
            12'd3977: current_page <= 12'd4095;
            12'd3978: current_page <= 12'd4095;
            12'd3979: current_page <= 12'd4095;
            12'd3980: current_page <= 12'd4095;
            12'd3981: current_page <= 12'd4095;
            12'd3982: current_page <= 12'd4095;
            12'd3983: current_page <= 12'd4095;
            12'd3984: current_page <= 12'd4095;
            12'd3985: current_page <= 12'd4095;
            12'd3986: current_page <= 12'd4095;
            12'd3987: current_page <= 12'd4095;
            12'd3988: current_page <= 12'd4095;
            12'd3989: current_page <= 12'd4095;
            12'd3990: current_page <= 12'd4095;
            12'd3991: current_page <= 12'd4095;
            12'd3992: current_page <= 12'd4095;
            12'd3993: current_page <= 12'd4095;
            12'd3994: current_page <= 12'd4095;
            12'd3995: current_page <= 12'd4095;
            12'd3996: current_page <= 12'd4095;
            12'd3997: current_page <= 12'd4095;
            12'd3998: current_page <= 12'd4095;
            12'd3999: current_page <= 12'd4095;
            12'd4000: current_page <= 12'd4095;
            12'd4001: current_page <= 12'd4095;
            12'd4002: current_page <= 12'd4095;
            12'd4003: current_page <= 12'd4095;
            12'd4004: current_page <= 12'd4095;
            12'd4005: current_page <= 12'd4095;
            12'd4006: current_page <= 12'd4095;
            12'd4007: current_page <= 12'd4095;
            12'd4008: current_page <= 12'd4095;
            12'd4009: current_page <= 12'd4095;
            12'd4010: current_page <= 12'd4095;
            12'd4011: current_page <= 12'd4095;
            12'd4012: current_page <= 12'd4095;
            12'd4013: current_page <= 12'd4095;
            12'd4014: current_page <= 12'd4095;
            12'd4015: current_page <= 12'd4095;
            12'd4016: current_page <= 12'd4095;
            12'd4017: current_page <= 12'd4095;
            12'd4018: current_page <= 12'd4095;
            12'd4019: current_page <= 12'd4095;
            12'd4020: current_page <= 12'd4095;
            12'd4021: current_page <= 12'd4095;
            12'd4022: current_page <= 12'd4095;
            12'd4023: current_page <= 12'd4095;
            12'd4024: current_page <= 12'd4095;
            12'd4025: current_page <= 12'd4095;
            12'd4026: current_page <= 12'd4095;
            12'd4027: current_page <= 12'd4095;
            12'd4028: current_page <= 12'd4095;
            12'd4029: current_page <= 12'd4095;
            12'd4030: current_page <= 12'd4095;
            12'd4031: current_page <= 12'd4095;
            12'd4032: current_page <= 12'd4095;
            12'd4033: current_page <= 12'd4095;
            12'd4034: current_page <= 12'd4095;
            12'd4035: current_page <= 12'd4095;
            12'd4036: current_page <= 12'd4095;
            12'd4037: current_page <= 12'd4095;
            12'd4038: current_page <= 12'd4095;
            12'd4039: current_page <= 12'd4095;
            12'd4040: current_page <= 12'd4095;
            12'd4041: current_page <= 12'd4095;
            12'd4042: current_page <= 12'd4095;
            12'd4043: current_page <= 12'd4095;
            12'd4044: current_page <= 12'd4095;
            12'd4045: current_page <= 12'd4095;
            12'd4046: current_page <= 12'd4095;
            12'd4047: current_page <= 12'd4095;
            12'd4048: current_page <= 12'd4095;
            12'd4049: current_page <= 12'd4095;
            12'd4050: current_page <= 12'd4095;
            12'd4051: current_page <= 12'd4095;
            12'd4052: current_page <= 12'd4095;
            12'd4053: current_page <= 12'd4095;
            12'd4054: current_page <= 12'd4095;
            12'd4055: current_page <= 12'd4095;
            12'd4056: current_page <= 12'd4095;
            12'd4057: current_page <= 12'd4095;
            12'd4058: current_page <= 12'd4095;
            12'd4059: current_page <= 12'd4095;
            12'd4060: current_page <= 12'd4095;
            12'd4061: current_page <= 12'd4095;
            12'd4062: current_page <= 12'd4095;
            12'd4063: current_page <= 12'd4095;
            12'd4064: current_page <= 12'd4095;
            12'd4065: current_page <= 12'd4095;
            12'd4066: current_page <= 12'd4095;
            12'd4067: current_page <= 12'd4095;
            12'd4068: current_page <= 12'd4095;
            12'd4069: current_page <= 12'd4095;
            12'd4070: current_page <= 12'd4095;
            12'd4071: current_page <= 12'd4095;
            12'd4072: current_page <= 12'd4095;
            12'd4073: current_page <= 12'd4095;
            12'd4074: current_page <= 12'd4095;
            12'd4075: current_page <= 12'd4095;
            12'd4076: current_page <= 12'd4095;
            12'd4077: current_page <= 12'd4095;
            12'd4078: current_page <= 12'd4095;
            12'd4079: current_page <= 12'd4095;
            12'd4080: current_page <= 12'd4095;
            12'd4081: current_page <= 12'd4095;
            12'd4082: current_page <= 12'd4095;
            12'd4083: current_page <= 12'd4095;
            12'd4084: current_page <= 12'd4095;
            12'd4085: current_page <= 12'd4095;
            12'd4086: current_page <= 12'd4095;
            12'd4087: current_page <= 12'd4095;
            12'd4088: current_page <= 12'd4095;
            12'd4089: current_page <= 12'd4095;
            12'd4090: current_page <= 12'd4095;
            12'd4091: current_page <= 12'd4095;
            12'd4092: current_page <= 12'd4095;
            12'd4093: current_page <= 12'd4095;
            12'd4094: current_page <= 12'd4095;
            12'd4095: current_page <= 12'd4095;
        endcase
    end
endmodule
